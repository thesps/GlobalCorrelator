../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/reduce_17.vhd