../../../../../../RuflCore/firmware/hdl/ReuseableElements/DataPipe.vhd