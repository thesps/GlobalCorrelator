../../../../../../HGC-firmware/projects/Common/firmware/hdl/ReuseableElements/PkgArrayTypes.vhd