../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/reduce_7.vhd