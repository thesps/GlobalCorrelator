../../../../../../../GlobalCorrelator_HLS/JetLoop/solution1/syn/vhdl/reduce_1.vhd