../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/jet_compute_mul_mdEe.vhd