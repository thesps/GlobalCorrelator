../../../../../../../RuflCore/firmware/hdl/ReuseableElements/DataRam.vhd