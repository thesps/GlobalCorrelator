../../../../../../HGC-firmware/projects/Common/firmware/hdl/ReuseableElements/DataPipe.vhd