library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library Utilities;
use Utilities.Utilities.all;

library Layer2;
use Layer2.Constants.all;

library PFChargedObj;
use PFChargedObj.DataType;
use PFChargedObj.ArrayTypes;

entity Seeding is
port(
  clk : in std_logic;
  PFChargedObjStream : in PFChargedObj.ArrayTypes.VectorPipe;
  Seeds : out PFChargedObj.ArrayTypes.VectorPipe
);
end Seeding;

architecture behavioral of Seeding is
  signal SeedsInt : PFChargedObj.ArrayTypes.Vector(0 to N_PF_Regions - 1) := PFChargedObj.ArrayTypes.NullVector(N_PF_Regions);
begin

-- Simplest, most naive seeding: take the highest pT object from each region
-- The objects arrive pT ordered so just take the first to arrvie
SeedGen:
--for i in 0 to N_PF_Regions - 1 generate
for i in 0 to N_PF_Regions_PerLayer1Board - 1 generate
begin
  process(clk)
  begin
  if rising_edge(clk) then
    if not PFChargedObjStream(1)(i).FrameValid and PFChargedObjStream(0)(i).FrameValid then
      SeedsInt(i) <= PFChargedObjStream(0)(i);
    end if;
  end if;
  end process;
end generate;

OutPipe : entity PFChargedObj.DataPipe
port map(clk, SeedsInt, Seeds);

DebugInstance : entity PFChargedObj.Debug
generic map( FileName => "Seeding" )
port map(clk, SeedsInt);

end behavioral;
