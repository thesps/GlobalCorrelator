library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library IO;
use IO.DataType.all;
use IO.ArrayTypes.all;

library JetLoop;

use work.PkgConstants.all;

entity JetLoopWrapped is
port(
    clk : in std_logic;
    particles_in : in Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    particles_out : out Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    in_cone : out Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    sum_pts : out Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    sum_pt_etas : out Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    sum_pt_phis : out Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    seed_eta : out tData := cNull;
    seed_phi : out tData := cNull
);
end JetLoopWrapped;

architecture rtl of JetLoopWrapped is

begin

    HLSIP : entity JetLoop.jet_loop
    port map(
    ap_clk => clk,
    ap_rst => '0',
    ap_start => '1',
    particles_in_0 => particles_in(0).data(35 downto 0),
    particles_in_1 => particles_in(1).data(35 downto 0),
    particles_in_2 => particles_in(2).data(35 downto 0),
    particles_in_3 => particles_in(3).data(35 downto 0),
    particles_in_4 => particles_in(4).data(35 downto 0),
    particles_in_5 => particles_in(5).data(35 downto 0),
    particles_in_6 => particles_in(6).data(35 downto 0),
    particles_in_7 => particles_in(7).data(35 downto 0),
    particles_in_8 => particles_in(8).data(35 downto 0),
    particles_in_9 => particles_in(9).data(35 downto 0),
    particles_in_10 => particles_in(10).data(35 downto 0),
    particles_in_11 => particles_in(11).data(35 downto 0),
    particles_in_12 => particles_in(12).data(35 downto 0),
    particles_in_13 => particles_in(13).data(35 downto 0),
    particles_in_14 => particles_in(14).data(35 downto 0),
    particles_in_15 => particles_in(15).data(35 downto 0),
    particles_in_16 => particles_in(16).data(35 downto 0),
    particles_in_17 => particles_in(17).data(35 downto 0),
    particles_in_18 => particles_in(18).data(35 downto 0),
    particles_in_19 => particles_in(19).data(35 downto 0),
    particles_in_20 => particles_in(20).data(35 downto 0),
    particles_in_21 => particles_in(21).data(35 downto 0),
    particles_in_22 => particles_in(22).data(35 downto 0),
    particles_in_23 => particles_in(23).data(35 downto 0),
    particles_in_24 => particles_in(24).data(35 downto 0),
    particles_in_25 => particles_in(25).data(35 downto 0),
    particles_in_26 => particles_in(26).data(35 downto 0),
    particles_in_27 => particles_in(27).data(35 downto 0),
    particles_in_28 => particles_in(28).data(35 downto 0),
    particles_in_29 => particles_in(29).data(35 downto 0),
    particles_in_30 => particles_in(30).data(35 downto 0),
    particles_in_31 => particles_in(31).data(35 downto 0),
    particles_in_32 => particles_in(32).data(35 downto 0),
    particles_in_33 => particles_in(33).data(35 downto 0),
    particles_in_34 => particles_in(34).data(35 downto 0),
    particles_in_35 => particles_in(35).data(35 downto 0),
    particles_in_36 => particles_in(36).data(35 downto 0),
    particles_in_37 => particles_in(37).data(35 downto 0),
    particles_in_38 => particles_in(38).data(35 downto 0),
    particles_in_39 => particles_in(39).data(35 downto 0),
    particles_in_40 => particles_in(40).data(35 downto 0),
    particles_in_41 => particles_in(41).data(35 downto 0),
    particles_in_42 => particles_in(42).data(35 downto 0),
    particles_in_43 => particles_in(43).data(35 downto 0),
    particles_in_44 => particles_in(44).data(35 downto 0),
    particles_in_45 => particles_in(45).data(35 downto 0),
    particles_in_46 => particles_in(46).data(35 downto 0),
    particles_in_47 => particles_in(47).data(35 downto 0),
    particles_in_48 => particles_in(48).data(35 downto 0),
    particles_in_49 => particles_in(49).data(35 downto 0),
    particles_in_50 => particles_in(50).data(35 downto 0),
    particles_in_51 => particles_in(51).data(35 downto 0),
    particles_in_52 => particles_in(52).data(35 downto 0),
    particles_in_53 => particles_in(53).data(35 downto 0),
    particles_in_54 => particles_in(54).data(35 downto 0),
    particles_in_55 => particles_in(55).data(35 downto 0),
    particles_in_56 => particles_in(56).data(35 downto 0),
    particles_in_57 => particles_in(57).data(35 downto 0),
    particles_in_58 => particles_in(58).data(35 downto 0),
    particles_in_59 => particles_in(59).data(35 downto 0),
    particles_in_60 => particles_in(60).data(35 downto 0),
    particles_in_61 => particles_in(61).data(35 downto 0),
    particles_in_62 => particles_in(62).data(35 downto 0),
    particles_in_63 => particles_in(63).data(35 downto 0),
    particles_in_64 => particles_in(64).data(35 downto 0),
    particles_in_65 => particles_in(65).data(35 downto 0),
    particles_in_66 => particles_in(66).data(35 downto 0),
    particles_in_67 => particles_in(67).data(35 downto 0),
    particles_in_68 => particles_in(68).data(35 downto 0),
    particles_in_69 => particles_in(69).data(35 downto 0),
    particles_in_70 => particles_in(70).data(35 downto 0),
    particles_in_71 => particles_in(71).data(35 downto 0),
    particles_in_72 => particles_in(72).data(35 downto 0),
    particles_in_73 => particles_in(73).data(35 downto 0),
    particles_in_74 => particles_in(74).data(35 downto 0),
    particles_in_75 => particles_in(75).data(35 downto 0),
    particles_in_76 => particles_in(76).data(35 downto 0),
    particles_in_77 => particles_in(77).data(35 downto 0),
    particles_in_78 => particles_in(78).data(35 downto 0),
    particles_in_79 => particles_in(79).data(35 downto 0),
    particles_in_80 => particles_in(80).data(35 downto 0),
    particles_in_81 => particles_in(81).data(35 downto 0),
    particles_in_82 => particles_in(82).data(35 downto 0),
    particles_in_83 => particles_in(83).data(35 downto 0),
    particles_in_84 => particles_in(84).data(35 downto 0),
    particles_in_85 => particles_in(85).data(35 downto 0),
    particles_in_86 => particles_in(86).data(35 downto 0),
    particles_in_87 => particles_in(87).data(35 downto 0),
    particles_in_88 => particles_in(88).data(35 downto 0),
    particles_in_89 => particles_in(89).data(35 downto 0),
    particles_in_90 => particles_in(90).data(35 downto 0),
    particles_in_91 => particles_in(91).data(35 downto 0),
    particles_in_92 => particles_in(92).data(35 downto 0),
    particles_in_93 => particles_in(93).data(35 downto 0),
    particles_in_94 => particles_in(94).data(35 downto 0),
    particles_in_95 => particles_in(95).data(35 downto 0),
    particles_in_96 => particles_in(96).data(35 downto 0),
    particles_in_97 => particles_in(97).data(35 downto 0),
    particles_in_98 => particles_in(98).data(35 downto 0),
    particles_in_99 => particles_in(99).data(35 downto 0),
    particles_in_100 => particles_in(100).data(35 downto 0),
    particles_in_101 => particles_in(101).data(35 downto 0),
    particles_in_102 => particles_in(102).data(35 downto 0),
    particles_in_103 => particles_in(103).data(35 downto 0),
    particles_in_104 => particles_in(104).data(35 downto 0),
    particles_in_105 => particles_in(105).data(35 downto 0),
    particles_in_106 => particles_in(106).data(35 downto 0),
    particles_in_107 => particles_in(107).data(35 downto 0),
    particles_in_108 => particles_in(108).data(35 downto 0),
    particles_in_109 => particles_in(109).data(35 downto 0),
    particles_in_110 => particles_in(110).data(35 downto 0),
    particles_in_111 => particles_in(111).data(35 downto 0),
    particles_in_112 => particles_in(112).data(35 downto 0),
    particles_in_113 => particles_in(113).data(35 downto 0),
    particles_in_114 => particles_in(114).data(35 downto 0),
    particles_in_115 => particles_in(115).data(35 downto 0),
    particles_in_116 => particles_in(116).data(35 downto 0),
    particles_in_117 => particles_in(117).data(35 downto 0),
    particles_in_118 => particles_in(118).data(35 downto 0),
    particles_in_119 => particles_in(119).data(35 downto 0),
    particles_in_120 => particles_in(120).data(35 downto 0),
    particles_in_121 => particles_in(121).data(35 downto 0),
    particles_in_122 => particles_in(122).data(35 downto 0),
    particles_in_123 => particles_in(123).data(35 downto 0),
    particles_in_124 => particles_in(124).data(35 downto 0),
    particles_in_125 => particles_in(125).data(35 downto 0),
    particles_in_126 => particles_in(126).data(35 downto 0),
    particles_in_127 => particles_in(127).data(35 downto 0),
    particles_out_0 => particles_out(0).data(35 downto 0),
    particles_out_1 => particles_out(1).data(35 downto 0),
    particles_out_2 => particles_out(2).data(35 downto 0),
    particles_out_3 => particles_out(3).data(35 downto 0),
    particles_out_4 => particles_out(4).data(35 downto 0),
    particles_out_5 => particles_out(5).data(35 downto 0),
    particles_out_6 => particles_out(6).data(35 downto 0),
    particles_out_7 => particles_out(7).data(35 downto 0),
    particles_out_8 => particles_out(8).data(35 downto 0),
    particles_out_9 => particles_out(9).data(35 downto 0),
    particles_out_10 => particles_out(10).data(35 downto 0),
    particles_out_11 => particles_out(11).data(35 downto 0),
    particles_out_12 => particles_out(12).data(35 downto 0),
    particles_out_13 => particles_out(13).data(35 downto 0),
    particles_out_14 => particles_out(14).data(35 downto 0),
    particles_out_15 => particles_out(15).data(35 downto 0),
    particles_out_16 => particles_out(16).data(35 downto 0),
    particles_out_17 => particles_out(17).data(35 downto 0),
    particles_out_18 => particles_out(18).data(35 downto 0),
    particles_out_19 => particles_out(19).data(35 downto 0),
    particles_out_20 => particles_out(20).data(35 downto 0),
    particles_out_21 => particles_out(21).data(35 downto 0),
    particles_out_22 => particles_out(22).data(35 downto 0),
    particles_out_23 => particles_out(23).data(35 downto 0),
    particles_out_24 => particles_out(24).data(35 downto 0),
    particles_out_25 => particles_out(25).data(35 downto 0),
    particles_out_26 => particles_out(26).data(35 downto 0),
    particles_out_27 => particles_out(27).data(35 downto 0),
    particles_out_28 => particles_out(28).data(35 downto 0),
    particles_out_29 => particles_out(29).data(35 downto 0),
    particles_out_30 => particles_out(30).data(35 downto 0),
    particles_out_31 => particles_out(31).data(35 downto 0),
    particles_out_32 => particles_out(32).data(35 downto 0),
    particles_out_33 => particles_out(33).data(35 downto 0),
    particles_out_34 => particles_out(34).data(35 downto 0),
    particles_out_35 => particles_out(35).data(35 downto 0),
    particles_out_36 => particles_out(36).data(35 downto 0),
    particles_out_37 => particles_out(37).data(35 downto 0),
    particles_out_38 => particles_out(38).data(35 downto 0),
    particles_out_39 => particles_out(39).data(35 downto 0),
    particles_out_40 => particles_out(40).data(35 downto 0),
    particles_out_41 => particles_out(41).data(35 downto 0),
    particles_out_42 => particles_out(42).data(35 downto 0),
    particles_out_43 => particles_out(43).data(35 downto 0),
    particles_out_44 => particles_out(44).data(35 downto 0),
    particles_out_45 => particles_out(45).data(35 downto 0),
    particles_out_46 => particles_out(46).data(35 downto 0),
    particles_out_47 => particles_out(47).data(35 downto 0),
    particles_out_48 => particles_out(48).data(35 downto 0),
    particles_out_49 => particles_out(49).data(35 downto 0),
    particles_out_50 => particles_out(50).data(35 downto 0),
    particles_out_51 => particles_out(51).data(35 downto 0),
    particles_out_52 => particles_out(52).data(35 downto 0),
    particles_out_53 => particles_out(53).data(35 downto 0),
    particles_out_54 => particles_out(54).data(35 downto 0),
    particles_out_55 => particles_out(55).data(35 downto 0),
    particles_out_56 => particles_out(56).data(35 downto 0),
    particles_out_57 => particles_out(57).data(35 downto 0),
    particles_out_58 => particles_out(58).data(35 downto 0),
    particles_out_59 => particles_out(59).data(35 downto 0),
    particles_out_60 => particles_out(60).data(35 downto 0),
    particles_out_61 => particles_out(61).data(35 downto 0),
    particles_out_62 => particles_out(62).data(35 downto 0),
    particles_out_63 => particles_out(63).data(35 downto 0),
    particles_out_64 => particles_out(64).data(35 downto 0),
    particles_out_65 => particles_out(65).data(35 downto 0),
    particles_out_66 => particles_out(66).data(35 downto 0),
    particles_out_67 => particles_out(67).data(35 downto 0),
    particles_out_68 => particles_out(68).data(35 downto 0),
    particles_out_69 => particles_out(69).data(35 downto 0),
    particles_out_70 => particles_out(70).data(35 downto 0),
    particles_out_71 => particles_out(71).data(35 downto 0),
    particles_out_72 => particles_out(72).data(35 downto 0),
    particles_out_73 => particles_out(73).data(35 downto 0),
    particles_out_74 => particles_out(74).data(35 downto 0),
    particles_out_75 => particles_out(75).data(35 downto 0),
    particles_out_76 => particles_out(76).data(35 downto 0),
    particles_out_77 => particles_out(77).data(35 downto 0),
    particles_out_78 => particles_out(78).data(35 downto 0),
    particles_out_79 => particles_out(79).data(35 downto 0),
    particles_out_80 => particles_out(80).data(35 downto 0),
    particles_out_81 => particles_out(81).data(35 downto 0),
    particles_out_82 => particles_out(82).data(35 downto 0),
    particles_out_83 => particles_out(83).data(35 downto 0),
    particles_out_84 => particles_out(84).data(35 downto 0),
    particles_out_85 => particles_out(85).data(35 downto 0),
    particles_out_86 => particles_out(86).data(35 downto 0),
    particles_out_87 => particles_out(87).data(35 downto 0),
    particles_out_88 => particles_out(88).data(35 downto 0),
    particles_out_89 => particles_out(89).data(35 downto 0),
    particles_out_90 => particles_out(90).data(35 downto 0),
    particles_out_91 => particles_out(91).data(35 downto 0),
    particles_out_92 => particles_out(92).data(35 downto 0),
    particles_out_93 => particles_out(93).data(35 downto 0),
    particles_out_94 => particles_out(94).data(35 downto 0),
    particles_out_95 => particles_out(95).data(35 downto 0),
    particles_out_96 => particles_out(96).data(35 downto 0),
    particles_out_97 => particles_out(97).data(35 downto 0),
    particles_out_98 => particles_out(98).data(35 downto 0),
    particles_out_99 => particles_out(99).data(35 downto 0),
    particles_out_100 => particles_out(100).data(35 downto 0),
    particles_out_101 => particles_out(101).data(35 downto 0),
    particles_out_102 => particles_out(102).data(35 downto 0),
    particles_out_103 => particles_out(103).data(35 downto 0),
    particles_out_104 => particles_out(104).data(35 downto 0),
    particles_out_105 => particles_out(105).data(35 downto 0),
    particles_out_106 => particles_out(106).data(35 downto 0),
    particles_out_107 => particles_out(107).data(35 downto 0),
    particles_out_108 => particles_out(108).data(35 downto 0),
    particles_out_109 => particles_out(109).data(35 downto 0),
    particles_out_110 => particles_out(110).data(35 downto 0),
    particles_out_111 => particles_out(111).data(35 downto 0),
    particles_out_112 => particles_out(112).data(35 downto 0),
    particles_out_113 => particles_out(113).data(35 downto 0),
    particles_out_114 => particles_out(114).data(35 downto 0),
    particles_out_115 => particles_out(115).data(35 downto 0),
    particles_out_116 => particles_out(116).data(35 downto 0),
    particles_out_117 => particles_out(117).data(35 downto 0),
    particles_out_118 => particles_out(118).data(35 downto 0),
    particles_out_119 => particles_out(119).data(35 downto 0),
    particles_out_120 => particles_out(120).data(35 downto 0),
    particles_out_121 => particles_out(121).data(35 downto 0),
    particles_out_122 => particles_out(122).data(35 downto 0),
    particles_out_123 => particles_out(123).data(35 downto 0),
    particles_out_124 => particles_out(124).data(35 downto 0),
    particles_out_125 => particles_out(125).data(35 downto 0),
    particles_out_126 => particles_out(126).data(35 downto 0),
    particles_out_127 => particles_out(127).data(35 downto 0),
    incone_0 => in_cone(0).data(0),
    incone_1 => in_cone(1).data(0),
    incone_2 => in_cone(2).data(0),
    incone_3 => in_cone(3).data(0),
    incone_4 => in_cone(4).data(0),
    incone_5 => in_cone(5).data(0),
    incone_6 => in_cone(6).data(0),
    incone_7 => in_cone(7).data(0),
    incone_8 => in_cone(8).data(0),
    incone_9 => in_cone(9).data(0),
    incone_10 => in_cone(10).data(0),
    incone_11 => in_cone(11).data(0),
    incone_12 => in_cone(12).data(0),
    incone_13 => in_cone(13).data(0),
    incone_14 => in_cone(14).data(0),
    incone_15 => in_cone(15).data(0),
    incone_16 => in_cone(16).data(0),
    incone_17 => in_cone(17).data(0),
    incone_18 => in_cone(18).data(0),
    incone_19 => in_cone(19).data(0),
    incone_20 => in_cone(20).data(0),
    incone_21 => in_cone(21).data(0),
    incone_22 => in_cone(22).data(0),
    incone_23 => in_cone(23).data(0),
    incone_24 => in_cone(24).data(0),
    incone_25 => in_cone(25).data(0),
    incone_26 => in_cone(26).data(0),
    incone_27 => in_cone(27).data(0),
    incone_28 => in_cone(28).data(0),
    incone_29 => in_cone(29).data(0),
    incone_30 => in_cone(30).data(0),
    incone_31 => in_cone(31).data(0),
    incone_32 => in_cone(32).data(0),
    incone_33 => in_cone(33).data(0),
    incone_34 => in_cone(34).data(0),
    incone_35 => in_cone(35).data(0),
    incone_36 => in_cone(36).data(0),
    incone_37 => in_cone(37).data(0),
    incone_38 => in_cone(38).data(0),
    incone_39 => in_cone(39).data(0),
    incone_40 => in_cone(40).data(0),
    incone_41 => in_cone(41).data(0),
    incone_42 => in_cone(42).data(0),
    incone_43 => in_cone(43).data(0),
    incone_44 => in_cone(44).data(0),
    incone_45 => in_cone(45).data(0),
    incone_46 => in_cone(46).data(0),
    incone_47 => in_cone(47).data(0),
    incone_48 => in_cone(48).data(0),
    incone_49 => in_cone(49).data(0),
    incone_50 => in_cone(50).data(0),
    incone_51 => in_cone(51).data(0),
    incone_52 => in_cone(52).data(0),
    incone_53 => in_cone(53).data(0),
    incone_54 => in_cone(54).data(0),
    incone_55 => in_cone(55).data(0),
    incone_56 => in_cone(56).data(0),
    incone_57 => in_cone(57).data(0),
    incone_58 => in_cone(58).data(0),
    incone_59 => in_cone(59).data(0),
    incone_60 => in_cone(60).data(0),
    incone_61 => in_cone(61).data(0),
    incone_62 => in_cone(62).data(0),
    incone_63 => in_cone(63).data(0),
    incone_64 => in_cone(64).data(0),
    incone_65 => in_cone(65).data(0),
    incone_66 => in_cone(66).data(0),
    incone_67 => in_cone(67).data(0),
    incone_68 => in_cone(68).data(0),
    incone_69 => in_cone(69).data(0),
    incone_70 => in_cone(70).data(0),
    incone_71 => in_cone(71).data(0),
    incone_72 => in_cone(72).data(0),
    incone_73 => in_cone(73).data(0),
    incone_74 => in_cone(74).data(0),
    incone_75 => in_cone(75).data(0),
    incone_76 => in_cone(76).data(0),
    incone_77 => in_cone(77).data(0),
    incone_78 => in_cone(78).data(0),
    incone_79 => in_cone(79).data(0),
    incone_80 => in_cone(80).data(0),
    incone_81 => in_cone(81).data(0),
    incone_82 => in_cone(82).data(0),
    incone_83 => in_cone(83).data(0),
    incone_84 => in_cone(84).data(0),
    incone_85 => in_cone(85).data(0),
    incone_86 => in_cone(86).data(0),
    incone_87 => in_cone(87).data(0),
    incone_88 => in_cone(88).data(0),
    incone_89 => in_cone(89).data(0),
    incone_90 => in_cone(90).data(0),
    incone_91 => in_cone(91).data(0),
    incone_92 => in_cone(92).data(0),
    incone_93 => in_cone(93).data(0),
    incone_94 => in_cone(94).data(0),
    incone_95 => in_cone(95).data(0),
    incone_96 => in_cone(96).data(0),
    incone_97 => in_cone(97).data(0),
    incone_98 => in_cone(98).data(0),
    incone_99 => in_cone(99).data(0),
    incone_100 => in_cone(100).data(0),
    incone_101 => in_cone(101).data(0),
    incone_102 => in_cone(102).data(0),
    incone_103 => in_cone(103).data(0),
    incone_104 => in_cone(104).data(0),
    incone_105 => in_cone(105).data(0),
    incone_106 => in_cone(106).data(0),
    incone_107 => in_cone(107).data(0),
    incone_108 => in_cone(108).data(0),
    incone_109 => in_cone(109).data(0),
    incone_110 => in_cone(110).data(0),
    incone_111 => in_cone(111).data(0),
    incone_112 => in_cone(112).data(0),
    incone_113 => in_cone(113).data(0),
    incone_114 => in_cone(114).data(0),
    incone_115 => in_cone(115).data(0),
    incone_116 => in_cone(116).data(0),
    incone_117 => in_cone(117).data(0),
    incone_118 => in_cone(118).data(0),
    incone_119 => in_cone(119).data(0),
    incone_120 => in_cone(120).data(0),
    incone_121 => in_cone(121).data(0),
    incone_122 => in_cone(122).data(0),
    incone_123 => in_cone(123).data(0),
    incone_124 => in_cone(124).data(0),
    incone_125 => in_cone(125).data(0),
    incone_126 => in_cone(126).data(0),
    incone_127 => in_cone(127).data(0),
    sum_pts_0_V => sum_pts(0).data(15 downto 0),
    sum_pts_1_V => sum_pts(1).data(15 downto 0),
    sum_pts_2_V => sum_pts(2).data(15 downto 0),
    sum_pts_3_V => sum_pts(3).data(15 downto 0),
    sum_pts_4_V => sum_pts(4).data(15 downto 0),
    sum_pts_5_V => sum_pts(5).data(15 downto 0),
    sum_pts_6_V => sum_pts(6).data(15 downto 0),
    sum_pts_7_V => sum_pts(7).data(15 downto 0),
    sum_pts_8_V => sum_pts(8).data(15 downto 0),
    sum_pts_9_V => sum_pts(9).data(15 downto 0),
    sum_pts_10_V => sum_pts(10).data(15 downto 0),
    sum_pts_11_V => sum_pts(11).data(15 downto 0),
    sum_pts_12_V => sum_pts(12).data(15 downto 0),
    sum_pts_13_V => sum_pts(13).data(15 downto 0),
    sum_pts_14_V => sum_pts(14).data(15 downto 0),
    sum_pts_15_V => sum_pts(15).data(15 downto 0),
    sum_pts_16_V => sum_pts(16).data(15 downto 0),
    sum_pts_17_V => sum_pts(17).data(15 downto 0),
    sum_pts_18_V => sum_pts(18).data(15 downto 0),
    sum_pts_19_V => sum_pts(19).data(15 downto 0),
    sum_pts_20_V => sum_pts(20).data(15 downto 0),
    sum_pts_21_V => sum_pts(21).data(15 downto 0),
    sum_pts_22_V => sum_pts(22).data(15 downto 0),
    sum_pts_23_V => sum_pts(23).data(15 downto 0),
    sum_pts_24_V => sum_pts(24).data(15 downto 0),
    sum_pts_25_V => sum_pts(25).data(15 downto 0),
    sum_pts_26_V => sum_pts(26).data(15 downto 0),
    sum_pts_27_V => sum_pts(27).data(15 downto 0),
    sum_pts_28_V => sum_pts(28).data(15 downto 0),
    sum_pts_29_V => sum_pts(29).data(15 downto 0),
    sum_pts_30_V => sum_pts(30).data(15 downto 0),
    sum_pts_31_V => sum_pts(31).data(15 downto 0),
    sum_pts_32_V => sum_pts(32).data(15 downto 0),
    sum_pts_33_V => sum_pts(33).data(15 downto 0),
    sum_pts_34_V => sum_pts(34).data(15 downto 0),
    sum_pts_35_V => sum_pts(35).data(15 downto 0),
    sum_pts_36_V => sum_pts(36).data(15 downto 0),
    sum_pts_37_V => sum_pts(37).data(15 downto 0),
    sum_pts_38_V => sum_pts(38).data(15 downto 0),
    sum_pts_39_V => sum_pts(39).data(15 downto 0),
    sum_pts_40_V => sum_pts(40).data(15 downto 0),
    sum_pts_41_V => sum_pts(41).data(15 downto 0),
    sum_pts_42_V => sum_pts(42).data(15 downto 0),
    sum_pts_43_V => sum_pts(43).data(15 downto 0),
    sum_pts_44_V => sum_pts(44).data(15 downto 0),
    sum_pts_45_V => sum_pts(45).data(15 downto 0),
    sum_pts_46_V => sum_pts(46).data(15 downto 0),
    sum_pts_47_V => sum_pts(47).data(15 downto 0),
    sum_pts_48_V => sum_pts(48).data(15 downto 0),
    sum_pts_49_V => sum_pts(49).data(15 downto 0),
    sum_pts_50_V => sum_pts(50).data(15 downto 0),
    sum_pts_51_V => sum_pts(51).data(15 downto 0),
    sum_pts_52_V => sum_pts(52).data(15 downto 0),
    sum_pts_53_V => sum_pts(53).data(15 downto 0),
    sum_pts_54_V => sum_pts(54).data(15 downto 0),
    sum_pts_55_V => sum_pts(55).data(15 downto 0),
    sum_pts_56_V => sum_pts(56).data(15 downto 0),
    sum_pts_57_V => sum_pts(57).data(15 downto 0),
    sum_pts_58_V => sum_pts(58).data(15 downto 0),
    sum_pts_59_V => sum_pts(59).data(15 downto 0),
    sum_pts_60_V => sum_pts(60).data(15 downto 0),
    sum_pts_61_V => sum_pts(61).data(15 downto 0),
    sum_pts_62_V => sum_pts(62).data(15 downto 0),
    sum_pts_63_V => sum_pts(63).data(15 downto 0),
    sum_pts_64_V => sum_pts(64).data(15 downto 0),
    sum_pts_65_V => sum_pts(65).data(15 downto 0),
    sum_pts_66_V => sum_pts(66).data(15 downto 0),
    sum_pts_67_V => sum_pts(67).data(15 downto 0),
    sum_pts_68_V => sum_pts(68).data(15 downto 0),
    sum_pts_69_V => sum_pts(69).data(15 downto 0),
    sum_pts_70_V => sum_pts(70).data(15 downto 0),
    sum_pts_71_V => sum_pts(71).data(15 downto 0),
    sum_pts_72_V => sum_pts(72).data(15 downto 0),
    sum_pts_73_V => sum_pts(73).data(15 downto 0),
    sum_pts_74_V => sum_pts(74).data(15 downto 0),
    sum_pts_75_V => sum_pts(75).data(15 downto 0),
    sum_pts_76_V => sum_pts(76).data(15 downto 0),
    sum_pts_77_V => sum_pts(77).data(15 downto 0),
    sum_pts_78_V => sum_pts(78).data(15 downto 0),
    sum_pts_79_V => sum_pts(79).data(15 downto 0),
    sum_pts_80_V => sum_pts(80).data(15 downto 0),
    sum_pts_81_V => sum_pts(81).data(15 downto 0),
    sum_pts_82_V => sum_pts(82).data(15 downto 0),
    sum_pts_83_V => sum_pts(83).data(15 downto 0),
    sum_pts_84_V => sum_pts(84).data(15 downto 0),
    sum_pts_85_V => sum_pts(85).data(15 downto 0),
    sum_pts_86_V => sum_pts(86).data(15 downto 0),
    sum_pts_87_V => sum_pts(87).data(15 downto 0),
    sum_pts_88_V => sum_pts(88).data(15 downto 0),
    sum_pts_89_V => sum_pts(89).data(15 downto 0),
    sum_pts_90_V => sum_pts(90).data(15 downto 0),
    sum_pts_91_V => sum_pts(91).data(15 downto 0),
    sum_pts_92_V => sum_pts(92).data(15 downto 0),
    sum_pts_93_V => sum_pts(93).data(15 downto 0),
    sum_pts_94_V => sum_pts(94).data(15 downto 0),
    sum_pts_95_V => sum_pts(95).data(15 downto 0),
    sum_pts_96_V => sum_pts(96).data(15 downto 0),
    sum_pts_97_V => sum_pts(97).data(15 downto 0),
    sum_pts_98_V => sum_pts(98).data(15 downto 0),
    sum_pts_99_V => sum_pts(99).data(15 downto 0),
    sum_pts_100_V => sum_pts(100).data(15 downto 0),
    sum_pts_101_V => sum_pts(101).data(15 downto 0),
    sum_pts_102_V => sum_pts(102).data(15 downto 0),
    sum_pts_103_V => sum_pts(103).data(15 downto 0),
    sum_pts_104_V => sum_pts(104).data(15 downto 0),
    sum_pts_105_V => sum_pts(105).data(15 downto 0),
    sum_pts_106_V => sum_pts(106).data(15 downto 0),
    sum_pts_107_V => sum_pts(107).data(15 downto 0),
    sum_pts_108_V => sum_pts(108).data(15 downto 0),
    sum_pts_109_V => sum_pts(109).data(15 downto 0),
    sum_pts_110_V => sum_pts(110).data(15 downto 0),
    sum_pts_111_V => sum_pts(111).data(15 downto 0),
    sum_pts_112_V => sum_pts(112).data(15 downto 0),
    sum_pts_113_V => sum_pts(113).data(15 downto 0),
    sum_pts_114_V => sum_pts(114).data(15 downto 0),
    sum_pts_115_V => sum_pts(115).data(15 downto 0),
    sum_pts_116_V => sum_pts(116).data(15 downto 0),
    sum_pts_117_V => sum_pts(117).data(15 downto 0),
    sum_pts_118_V => sum_pts(118).data(15 downto 0),
    sum_pts_119_V => sum_pts(119).data(15 downto 0),
    sum_pts_120_V => sum_pts(120).data(15 downto 0),
    sum_pts_121_V => sum_pts(121).data(15 downto 0),
    sum_pts_122_V => sum_pts(122).data(15 downto 0),
    sum_pts_123_V => sum_pts(123).data(15 downto 0),
    sum_pts_124_V => sum_pts(124).data(15 downto 0),
    sum_pts_125_V => sum_pts(125).data(15 downto 0),
    sum_pts_126_V => sum_pts(126).data(15 downto 0),
    sum_pts_127_V => sum_pts(127).data(15 downto 0),
    sum_pt_etas_0_V => sum_pt_etas(0).data(21 downto 0),
    sum_pt_etas_1_V => sum_pt_etas(1).data(21 downto 0),
    sum_pt_etas_2_V => sum_pt_etas(2).data(21 downto 0),
    sum_pt_etas_3_V => sum_pt_etas(3).data(21 downto 0),
    sum_pt_etas_4_V => sum_pt_etas(4).data(21 downto 0),
    sum_pt_etas_5_V => sum_pt_etas(5).data(21 downto 0),
    sum_pt_etas_6_V => sum_pt_etas(6).data(21 downto 0),
    sum_pt_etas_7_V => sum_pt_etas(7).data(21 downto 0),
    sum_pt_etas_8_V => sum_pt_etas(8).data(21 downto 0),
    sum_pt_etas_9_V => sum_pt_etas(9).data(21 downto 0),
    sum_pt_etas_10_V => sum_pt_etas(10).data(21 downto 0),
    sum_pt_etas_11_V => sum_pt_etas(11).data(21 downto 0),
    sum_pt_etas_12_V => sum_pt_etas(12).data(21 downto 0),
    sum_pt_etas_13_V => sum_pt_etas(13).data(21 downto 0),
    sum_pt_etas_14_V => sum_pt_etas(14).data(21 downto 0),
    sum_pt_etas_15_V => sum_pt_etas(15).data(21 downto 0),
    sum_pt_etas_16_V => sum_pt_etas(16).data(21 downto 0),
    sum_pt_etas_17_V => sum_pt_etas(17).data(21 downto 0),
    sum_pt_etas_18_V => sum_pt_etas(18).data(21 downto 0),
    sum_pt_etas_19_V => sum_pt_etas(19).data(21 downto 0),
    sum_pt_etas_20_V => sum_pt_etas(20).data(21 downto 0),
    sum_pt_etas_21_V => sum_pt_etas(21).data(21 downto 0),
    sum_pt_etas_22_V => sum_pt_etas(22).data(21 downto 0),
    sum_pt_etas_23_V => sum_pt_etas(23).data(21 downto 0),
    sum_pt_etas_24_V => sum_pt_etas(24).data(21 downto 0),
    sum_pt_etas_25_V => sum_pt_etas(25).data(21 downto 0),
    sum_pt_etas_26_V => sum_pt_etas(26).data(21 downto 0),
    sum_pt_etas_27_V => sum_pt_etas(27).data(21 downto 0),
    sum_pt_etas_28_V => sum_pt_etas(28).data(21 downto 0),
    sum_pt_etas_29_V => sum_pt_etas(29).data(21 downto 0),
    sum_pt_etas_30_V => sum_pt_etas(30).data(21 downto 0),
    sum_pt_etas_31_V => sum_pt_etas(31).data(21 downto 0),
    sum_pt_etas_32_V => sum_pt_etas(32).data(21 downto 0),
    sum_pt_etas_33_V => sum_pt_etas(33).data(21 downto 0),
    sum_pt_etas_34_V => sum_pt_etas(34).data(21 downto 0),
    sum_pt_etas_35_V => sum_pt_etas(35).data(21 downto 0),
    sum_pt_etas_36_V => sum_pt_etas(36).data(21 downto 0),
    sum_pt_etas_37_V => sum_pt_etas(37).data(21 downto 0),
    sum_pt_etas_38_V => sum_pt_etas(38).data(21 downto 0),
    sum_pt_etas_39_V => sum_pt_etas(39).data(21 downto 0),
    sum_pt_etas_40_V => sum_pt_etas(40).data(21 downto 0),
    sum_pt_etas_41_V => sum_pt_etas(41).data(21 downto 0),
    sum_pt_etas_42_V => sum_pt_etas(42).data(21 downto 0),
    sum_pt_etas_43_V => sum_pt_etas(43).data(21 downto 0),
    sum_pt_etas_44_V => sum_pt_etas(44).data(21 downto 0),
    sum_pt_etas_45_V => sum_pt_etas(45).data(21 downto 0),
    sum_pt_etas_46_V => sum_pt_etas(46).data(21 downto 0),
    sum_pt_etas_47_V => sum_pt_etas(47).data(21 downto 0),
    sum_pt_etas_48_V => sum_pt_etas(48).data(21 downto 0),
    sum_pt_etas_49_V => sum_pt_etas(49).data(21 downto 0),
    sum_pt_etas_50_V => sum_pt_etas(50).data(21 downto 0),
    sum_pt_etas_51_V => sum_pt_etas(51).data(21 downto 0),
    sum_pt_etas_52_V => sum_pt_etas(52).data(21 downto 0),
    sum_pt_etas_53_V => sum_pt_etas(53).data(21 downto 0),
    sum_pt_etas_54_V => sum_pt_etas(54).data(21 downto 0),
    sum_pt_etas_55_V => sum_pt_etas(55).data(21 downto 0),
    sum_pt_etas_56_V => sum_pt_etas(56).data(21 downto 0),
    sum_pt_etas_57_V => sum_pt_etas(57).data(21 downto 0),
    sum_pt_etas_58_V => sum_pt_etas(58).data(21 downto 0),
    sum_pt_etas_59_V => sum_pt_etas(59).data(21 downto 0),
    sum_pt_etas_60_V => sum_pt_etas(60).data(21 downto 0),
    sum_pt_etas_61_V => sum_pt_etas(61).data(21 downto 0),
    sum_pt_etas_62_V => sum_pt_etas(62).data(21 downto 0),
    sum_pt_etas_63_V => sum_pt_etas(63).data(21 downto 0),
    sum_pt_etas_64_V => sum_pt_etas(64).data(21 downto 0),
    sum_pt_etas_65_V => sum_pt_etas(65).data(21 downto 0),
    sum_pt_etas_66_V => sum_pt_etas(66).data(21 downto 0),
    sum_pt_etas_67_V => sum_pt_etas(67).data(21 downto 0),
    sum_pt_etas_68_V => sum_pt_etas(68).data(21 downto 0),
    sum_pt_etas_69_V => sum_pt_etas(69).data(21 downto 0),
    sum_pt_etas_70_V => sum_pt_etas(70).data(21 downto 0),
    sum_pt_etas_71_V => sum_pt_etas(71).data(21 downto 0),
    sum_pt_etas_72_V => sum_pt_etas(72).data(21 downto 0),
    sum_pt_etas_73_V => sum_pt_etas(73).data(21 downto 0),
    sum_pt_etas_74_V => sum_pt_etas(74).data(21 downto 0),
    sum_pt_etas_75_V => sum_pt_etas(75).data(21 downto 0),
    sum_pt_etas_76_V => sum_pt_etas(76).data(21 downto 0),
    sum_pt_etas_77_V => sum_pt_etas(77).data(21 downto 0),
    sum_pt_etas_78_V => sum_pt_etas(78).data(21 downto 0),
    sum_pt_etas_79_V => sum_pt_etas(79).data(21 downto 0),
    sum_pt_etas_80_V => sum_pt_etas(80).data(21 downto 0),
    sum_pt_etas_81_V => sum_pt_etas(81).data(21 downto 0),
    sum_pt_etas_82_V => sum_pt_etas(82).data(21 downto 0),
    sum_pt_etas_83_V => sum_pt_etas(83).data(21 downto 0),
    sum_pt_etas_84_V => sum_pt_etas(84).data(21 downto 0),
    sum_pt_etas_85_V => sum_pt_etas(85).data(21 downto 0),
    sum_pt_etas_86_V => sum_pt_etas(86).data(21 downto 0),
    sum_pt_etas_87_V => sum_pt_etas(87).data(21 downto 0),
    sum_pt_etas_88_V => sum_pt_etas(88).data(21 downto 0),
    sum_pt_etas_89_V => sum_pt_etas(89).data(21 downto 0),
    sum_pt_etas_90_V => sum_pt_etas(90).data(21 downto 0),
    sum_pt_etas_91_V => sum_pt_etas(91).data(21 downto 0),
    sum_pt_etas_92_V => sum_pt_etas(92).data(21 downto 0),
    sum_pt_etas_93_V => sum_pt_etas(93).data(21 downto 0),
    sum_pt_etas_94_V => sum_pt_etas(94).data(21 downto 0),
    sum_pt_etas_95_V => sum_pt_etas(95).data(21 downto 0),
    sum_pt_etas_96_V => sum_pt_etas(96).data(21 downto 0),
    sum_pt_etas_97_V => sum_pt_etas(97).data(21 downto 0),
    sum_pt_etas_98_V => sum_pt_etas(98).data(21 downto 0),
    sum_pt_etas_99_V => sum_pt_etas(99).data(21 downto 0),
    sum_pt_etas_100_V => sum_pt_etas(100).data(21 downto 0),
    sum_pt_etas_101_V => sum_pt_etas(101).data(21 downto 0),
    sum_pt_etas_102_V => sum_pt_etas(102).data(21 downto 0),
    sum_pt_etas_103_V => sum_pt_etas(103).data(21 downto 0),
    sum_pt_etas_104_V => sum_pt_etas(104).data(21 downto 0),
    sum_pt_etas_105_V => sum_pt_etas(105).data(21 downto 0),
    sum_pt_etas_106_V => sum_pt_etas(106).data(21 downto 0),
    sum_pt_etas_107_V => sum_pt_etas(107).data(21 downto 0),
    sum_pt_etas_108_V => sum_pt_etas(108).data(21 downto 0),
    sum_pt_etas_109_V => sum_pt_etas(109).data(21 downto 0),
    sum_pt_etas_110_V => sum_pt_etas(110).data(21 downto 0),
    sum_pt_etas_111_V => sum_pt_etas(111).data(21 downto 0),
    sum_pt_etas_112_V => sum_pt_etas(112).data(21 downto 0),
    sum_pt_etas_113_V => sum_pt_etas(113).data(21 downto 0),
    sum_pt_etas_114_V => sum_pt_etas(114).data(21 downto 0),
    sum_pt_etas_115_V => sum_pt_etas(115).data(21 downto 0),
    sum_pt_etas_116_V => sum_pt_etas(116).data(21 downto 0),
    sum_pt_etas_117_V => sum_pt_etas(117).data(21 downto 0),
    sum_pt_etas_118_V => sum_pt_etas(118).data(21 downto 0),
    sum_pt_etas_119_V => sum_pt_etas(119).data(21 downto 0),
    sum_pt_etas_120_V => sum_pt_etas(120).data(21 downto 0),
    sum_pt_etas_121_V => sum_pt_etas(121).data(21 downto 0),
    sum_pt_etas_122_V => sum_pt_etas(122).data(21 downto 0),
    sum_pt_etas_123_V => sum_pt_etas(123).data(21 downto 0),
    sum_pt_etas_124_V => sum_pt_etas(124).data(21 downto 0),
    sum_pt_etas_125_V => sum_pt_etas(125).data(21 downto 0),
    sum_pt_etas_126_V => sum_pt_etas(126).data(21 downto 0),
    sum_pt_etas_127_V => sum_pt_etas(127).data(21 downto 0),
    sum_pt_phis_0_V => sum_pt_phis(0).data(21 downto 0),
    sum_pt_phis_1_V => sum_pt_phis(1).data(21 downto 0),
    sum_pt_phis_2_V => sum_pt_phis(2).data(21 downto 0),
    sum_pt_phis_3_V => sum_pt_phis(3).data(21 downto 0),
    sum_pt_phis_4_V => sum_pt_phis(4).data(21 downto 0),
    sum_pt_phis_5_V => sum_pt_phis(5).data(21 downto 0),
    sum_pt_phis_6_V => sum_pt_phis(6).data(21 downto 0),
    sum_pt_phis_7_V => sum_pt_phis(7).data(21 downto 0),
    sum_pt_phis_8_V => sum_pt_phis(8).data(21 downto 0),
    sum_pt_phis_9_V => sum_pt_phis(9).data(21 downto 0),
    sum_pt_phis_10_V => sum_pt_phis(10).data(21 downto 0),
    sum_pt_phis_11_V => sum_pt_phis(11).data(21 downto 0),
    sum_pt_phis_12_V => sum_pt_phis(12).data(21 downto 0),
    sum_pt_phis_13_V => sum_pt_phis(13).data(21 downto 0),
    sum_pt_phis_14_V => sum_pt_phis(14).data(21 downto 0),
    sum_pt_phis_15_V => sum_pt_phis(15).data(21 downto 0),
    sum_pt_phis_16_V => sum_pt_phis(16).data(21 downto 0),
    sum_pt_phis_17_V => sum_pt_phis(17).data(21 downto 0),
    sum_pt_phis_18_V => sum_pt_phis(18).data(21 downto 0),
    sum_pt_phis_19_V => sum_pt_phis(19).data(21 downto 0),
    sum_pt_phis_20_V => sum_pt_phis(20).data(21 downto 0),
    sum_pt_phis_21_V => sum_pt_phis(21).data(21 downto 0),
    sum_pt_phis_22_V => sum_pt_phis(22).data(21 downto 0),
    sum_pt_phis_23_V => sum_pt_phis(23).data(21 downto 0),
    sum_pt_phis_24_V => sum_pt_phis(24).data(21 downto 0),
    sum_pt_phis_25_V => sum_pt_phis(25).data(21 downto 0),
    sum_pt_phis_26_V => sum_pt_phis(26).data(21 downto 0),
    sum_pt_phis_27_V => sum_pt_phis(27).data(21 downto 0),
    sum_pt_phis_28_V => sum_pt_phis(28).data(21 downto 0),
    sum_pt_phis_29_V => sum_pt_phis(29).data(21 downto 0),
    sum_pt_phis_30_V => sum_pt_phis(30).data(21 downto 0),
    sum_pt_phis_31_V => sum_pt_phis(31).data(21 downto 0),
    sum_pt_phis_32_V => sum_pt_phis(32).data(21 downto 0),
    sum_pt_phis_33_V => sum_pt_phis(33).data(21 downto 0),
    sum_pt_phis_34_V => sum_pt_phis(34).data(21 downto 0),
    sum_pt_phis_35_V => sum_pt_phis(35).data(21 downto 0),
    sum_pt_phis_36_V => sum_pt_phis(36).data(21 downto 0),
    sum_pt_phis_37_V => sum_pt_phis(37).data(21 downto 0),
    sum_pt_phis_38_V => sum_pt_phis(38).data(21 downto 0),
    sum_pt_phis_39_V => sum_pt_phis(39).data(21 downto 0),
    sum_pt_phis_40_V => sum_pt_phis(40).data(21 downto 0),
    sum_pt_phis_41_V => sum_pt_phis(41).data(21 downto 0),
    sum_pt_phis_42_V => sum_pt_phis(42).data(21 downto 0),
    sum_pt_phis_43_V => sum_pt_phis(43).data(21 downto 0),
    sum_pt_phis_44_V => sum_pt_phis(44).data(21 downto 0),
    sum_pt_phis_45_V => sum_pt_phis(45).data(21 downto 0),
    sum_pt_phis_46_V => sum_pt_phis(46).data(21 downto 0),
    sum_pt_phis_47_V => sum_pt_phis(47).data(21 downto 0),
    sum_pt_phis_48_V => sum_pt_phis(48).data(21 downto 0),
    sum_pt_phis_49_V => sum_pt_phis(49).data(21 downto 0),
    sum_pt_phis_50_V => sum_pt_phis(50).data(21 downto 0),
    sum_pt_phis_51_V => sum_pt_phis(51).data(21 downto 0),
    sum_pt_phis_52_V => sum_pt_phis(52).data(21 downto 0),
    sum_pt_phis_53_V => sum_pt_phis(53).data(21 downto 0),
    sum_pt_phis_54_V => sum_pt_phis(54).data(21 downto 0),
    sum_pt_phis_55_V => sum_pt_phis(55).data(21 downto 0),
    sum_pt_phis_56_V => sum_pt_phis(56).data(21 downto 0),
    sum_pt_phis_57_V => sum_pt_phis(57).data(21 downto 0),
    sum_pt_phis_58_V => sum_pt_phis(58).data(21 downto 0),
    sum_pt_phis_59_V => sum_pt_phis(59).data(21 downto 0),
    sum_pt_phis_60_V => sum_pt_phis(60).data(21 downto 0),
    sum_pt_phis_61_V => sum_pt_phis(61).data(21 downto 0),
    sum_pt_phis_62_V => sum_pt_phis(62).data(21 downto 0),
    sum_pt_phis_63_V => sum_pt_phis(63).data(21 downto 0),
    sum_pt_phis_64_V => sum_pt_phis(64).data(21 downto 0),
    sum_pt_phis_65_V => sum_pt_phis(65).data(21 downto 0),
    sum_pt_phis_66_V => sum_pt_phis(66).data(21 downto 0),
    sum_pt_phis_67_V => sum_pt_phis(67).data(21 downto 0),
    sum_pt_phis_68_V => sum_pt_phis(68).data(21 downto 0),
    sum_pt_phis_69_V => sum_pt_phis(69).data(21 downto 0),
    sum_pt_phis_70_V => sum_pt_phis(70).data(21 downto 0),
    sum_pt_phis_71_V => sum_pt_phis(71).data(21 downto 0),
    sum_pt_phis_72_V => sum_pt_phis(72).data(21 downto 0),
    sum_pt_phis_73_V => sum_pt_phis(73).data(21 downto 0),
    sum_pt_phis_74_V => sum_pt_phis(74).data(21 downto 0),
    sum_pt_phis_75_V => sum_pt_phis(75).data(21 downto 0),
    sum_pt_phis_76_V => sum_pt_phis(76).data(21 downto 0),
    sum_pt_phis_77_V => sum_pt_phis(77).data(21 downto 0),
    sum_pt_phis_78_V => sum_pt_phis(78).data(21 downto 0),
    sum_pt_phis_79_V => sum_pt_phis(79).data(21 downto 0),
    sum_pt_phis_80_V => sum_pt_phis(80).data(21 downto 0),
    sum_pt_phis_81_V => sum_pt_phis(81).data(21 downto 0),
    sum_pt_phis_82_V => sum_pt_phis(82).data(21 downto 0),
    sum_pt_phis_83_V => sum_pt_phis(83).data(21 downto 0),
    sum_pt_phis_84_V => sum_pt_phis(84).data(21 downto 0),
    sum_pt_phis_85_V => sum_pt_phis(85).data(21 downto 0),
    sum_pt_phis_86_V => sum_pt_phis(86).data(21 downto 0),
    sum_pt_phis_87_V => sum_pt_phis(87).data(21 downto 0),
    sum_pt_phis_88_V => sum_pt_phis(88).data(21 downto 0),
    sum_pt_phis_89_V => sum_pt_phis(89).data(21 downto 0),
    sum_pt_phis_90_V => sum_pt_phis(90).data(21 downto 0),
    sum_pt_phis_91_V => sum_pt_phis(91).data(21 downto 0),
    sum_pt_phis_92_V => sum_pt_phis(92).data(21 downto 0),
    sum_pt_phis_93_V => sum_pt_phis(93).data(21 downto 0),
    sum_pt_phis_94_V => sum_pt_phis(94).data(21 downto 0),
    sum_pt_phis_95_V => sum_pt_phis(95).data(21 downto 0),
    sum_pt_phis_96_V => sum_pt_phis(96).data(21 downto 0),
    sum_pt_phis_97_V => sum_pt_phis(97).data(21 downto 0),
    sum_pt_phis_98_V => sum_pt_phis(98).data(21 downto 0),
    sum_pt_phis_99_V => sum_pt_phis(99).data(21 downto 0),
    sum_pt_phis_100_V => sum_pt_phis(100).data(21 downto 0),
    sum_pt_phis_101_V => sum_pt_phis(101).data(21 downto 0),
    sum_pt_phis_102_V => sum_pt_phis(102).data(21 downto 0),
    sum_pt_phis_103_V => sum_pt_phis(103).data(21 downto 0),
    sum_pt_phis_104_V => sum_pt_phis(104).data(21 downto 0),
    sum_pt_phis_105_V => sum_pt_phis(105).data(21 downto 0),
    sum_pt_phis_106_V => sum_pt_phis(106).data(21 downto 0),
    sum_pt_phis_107_V => sum_pt_phis(107).data(21 downto 0),
    sum_pt_phis_108_V => sum_pt_phis(108).data(21 downto 0),
    sum_pt_phis_109_V => sum_pt_phis(109).data(21 downto 0),
    sum_pt_phis_110_V => sum_pt_phis(110).data(21 downto 0),
    sum_pt_phis_111_V => sum_pt_phis(111).data(21 downto 0),
    sum_pt_phis_112_V => sum_pt_phis(112).data(21 downto 0),
    sum_pt_phis_113_V => sum_pt_phis(113).data(21 downto 0),
    sum_pt_phis_114_V => sum_pt_phis(114).data(21 downto 0),
    sum_pt_phis_115_V => sum_pt_phis(115).data(21 downto 0),
    sum_pt_phis_116_V => sum_pt_phis(116).data(21 downto 0),
    sum_pt_phis_117_V => sum_pt_phis(117).data(21 downto 0),
    sum_pt_phis_118_V => sum_pt_phis(118).data(21 downto 0),
    sum_pt_phis_119_V => sum_pt_phis(119).data(21 downto 0),
    sum_pt_phis_120_V => sum_pt_phis(120).data(21 downto 0),
    sum_pt_phis_121_V => sum_pt_phis(121).data(21 downto 0),
    sum_pt_phis_122_V => sum_pt_phis(122).data(21 downto 0),
    sum_pt_phis_123_V => sum_pt_phis(123).data(21 downto 0),
    sum_pt_phis_124_V => sum_pt_phis(124).data(21 downto 0),
    sum_pt_phis_125_V => sum_pt_phis(125).data(21 downto 0),
    sum_pt_phis_126_V => sum_pt_phis(126).data(21 downto 0),
    sum_pt_phis_127_V => sum_pt_phis(127).data(21 downto 0),
    seed_eta_V => seed_eta.data(9 downto 0),
    seed_phi_V => seed_phi.data(9 downto 0)
    );

end rtl;
