library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Define constants related to the package
package PkgFindIndexInRow is

    constant moduleLatency : integer := 3;

end PkgFindIndexInRow;
