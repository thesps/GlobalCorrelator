../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/reduce_18.vhd