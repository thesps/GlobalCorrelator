../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/reduce_6.vhd