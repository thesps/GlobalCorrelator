../../../../../../../GlobalCorrelator_HLS/JetLoop/solution1/syn/vhdl/jet_loop.vhd