../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/reduce_19.vhd