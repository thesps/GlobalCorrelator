../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/jet_compute_inv_tbkb.vhd