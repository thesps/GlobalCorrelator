library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library Layer2;
use Layer2.Constants.all;

package Regions is

  -- Every region has 8 neighbours
  type NeighbourArray is array (0 to N_PF_Regions - 1, 0 to 8) of integer range -1 to N_PF_Regions - 1;
  constant Neighbours : NeighbourArray := 
((-1, -1, -1, 8, 0, 1, 17, 9, 10),
(-1, -1, -1, 0, 1, 2, 9, 10, 11),
(-1, -1, -1, 1, 2, 3, 10, 11, 12),
(-1, -1, -1, 2, 3, 4, 11, 12, 13),
(-1, -1, -1, 3, 4, 5, 12, 13, 14),
(-1, -1, -1, 4, 5, 6, 13, 14, 15),
(-1, -1, -1, 5, 6, 7, 14, 15, 16),
(-1, -1, -1, 6, 7, 8, 15, 16, 17),
(-1, -1, -1, 7, 8, 0, 16, 17, 9),
(8, 0, 1, 17, 9, 10, 26, 18, 19),
(0, 1, 2, 9, 10, 11, 18, 19, 20),
(1, 2, 3, 10, 11, 12, 19, 20, 21),
(2, 3, 4, 11, 12, 13, 20, 21, 22),
(3, 4, 5, 12, 13, 14, 21, 22, 23),
(4, 5, 6, 13, 14, 15, 22, 23, 24),
(5, 6, 7, 14, 15, 16, 23, 24, 25),
(6, 7, 8, 15, 16, 17, 24, 25, 26),
(7, 8, 0, 16, 17, 9, 25, 26, 18),
(17, 9, 10, 26, 18, 19, 35, 27, 28),
(9, 10, 11, 18, 19, 20, 27, 28, 29),
(10, 11, 12, 19, 20, 21, 28, 29, 30),
(11, 12, 13, 20, 21, 22, 29, 30, 31),
(12, 13, 14, 21, 22, 23, 30, 31, 32),
(13, 14, 15, 22, 23, 24, 31, 32, 33),
(14, 15, 16, 23, 24, 25, 32, 33, 34),
(15, 16, 17, 24, 25, 26, 33, 34, 35),
(16, 17, 9, 25, 26, 18, 34, 35, 27),
(26, 18, 19, 35, 27, 28, 44, 36, 37),
(18, 19, 20, 27, 28, 29, 36, 37, 38),
(19, 20, 21, 28, 29, 30, 37, 38, 39),
(20, 21, 22, 29, 30, 31, 38, 39, 40),
(21, 22, 23, 30, 31, 32, 39, 40, 41),
(22, 23, 24, 31, 32, 33, 40, 41, 42),
(23, 24, 25, 32, 33, 34, 41, 42, 43),
(24, 25, 26, 33, 34, 35, 42, 43, 44),
(25, 26, 18, 34, 35, 27, 43, 44, 36),
(35, 27, 28, 44, 36, 37, 53, 45, 46),
(27, 28, 29, 36, 37, 38, 45, 46, 47),
(28, 29, 30, 37, 38, 39, 46, 47, 48),
(29, 30, 31, 38, 39, 40, 47, 48, 49),
(30, 31, 32, 39, 40, 41, 48, 49, 50),
(31, 32, 33, 40, 41, 42, 49, 50, 51),
(32, 33, 34, 41, 42, 43, 50, 51, 52),
(33, 34, 35, 42, 43, 44, 51, 52, 53),
(34, 35, 27, 43, 44, 36, 52, 53, 45),
(44, 36, 37, 53, 45, 46, 62, 54, 55),
(36, 37, 38, 45, 46, 47, 54, 55, 56),
(37, 38, 39, 46, 47, 48, 55, 56, 57),
(38, 39, 40, 47, 48, 49, 56, 57, 58),
(39, 40, 41, 48, 49, 50, 57, 58, 59),
(40, 41, 42, 49, 50, 51, 58, 59, 60),
(41, 42, 43, 50, 51, 52, 59, 60, 61),
(42, 43, 44, 51, 52, 53, 60, 61, 62),
(43, 44, 36, 52, 53, 45, 61, 62, 54),
(53, 45, 46, 62, 54, 55, 71, 63, 64),
(45, 46, 47, 54, 55, 56, 63, 64, 65),
(46, 47, 48, 55, 56, 57, 64, 65, 66),
(47, 48, 49, 56, 57, 58, 65, 66, 67),
(48, 49, 50, 57, 58, 59, 66, 67, 68),
(49, 50, 51, 58, 59, 60, 67, 68, 69),
(50, 51, 52, 59, 60, 61, 68, 69, 70),
(51, 52, 53, 60, 61, 62, 69, 70, 71),
(52, 53, 45, 61, 62, 54, 70, 71, 63),
(62, 54, 55, 71, 63, 64, -1, -1, -1),
(54, 55, 56, 63, 64, 65, -1, -1, -1),
(55, 56, 57, 64, 65, 66, -1, -1, -1),
(56, 57, 58, 65, 66, 67, -1, -1, -1),
(57, 58, 59, 66, 67, 68, -1, -1, -1),
(58, 59, 60, 67, 68, 69, -1, -1, -1),
(59, 60, 61, 68, 69, 70, -1, -1, -1),
(60, 61, 62, 69, 70, 71, -1, -1, -1),
(61, 62, 54, 70, 71, 63, -1, -1, -1));

end Regions;
