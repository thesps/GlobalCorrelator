library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Constants is

    constant N_LINKS_HGC_TOTAL : integer := 12;
    constant N_REGIONS_PF : integer := 18;

end Constants;
