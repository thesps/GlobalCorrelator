../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/reduce_3.vhd