../../../../../../../GlobalCorrelator_HLS/JetCompute/solution1/syn/vhdl/jet_compute.vhd