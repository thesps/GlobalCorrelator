package pf_ip_constants is

  constant PF_ALGO_LATENCY : integer := 288;

end;
