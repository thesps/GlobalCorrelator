../../../../../../../RuflCore/firmware/hdl/ReuseableElements/Debugger.vhd