../../../../../../../GlobalCorrelator_HLS/JetLoop/solution1/syn/vhdl/reduce_2.vhd