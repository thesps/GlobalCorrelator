../../../../../../../GlobalCorrelator_HLS/JetLoop/solution1/syn/vhdl/reduce_6.vhd