../../../../../../../GlobalCorrelator_HLS/JetLoop/solution1/syn/vhdl/reduce_5.vhd