../../../../../../HGC-firmware/projects/Common/firmware/hdl/ReuseableElements/PairReduceMax.vhd