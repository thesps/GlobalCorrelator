library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pf_constants is

  constant PF_ALGO_LATENCY : natural := 91;  -- Algorithm latency in 240 MHz
                                             -- ticks
  --constant MAX_PF_IP_CORES : natural := 6;
  constant N_PF_IP_CORES : natural := 1;  -- Up to 6
  constant N_PF_IP_CORE_IN_CHANS : natural := 42;
  constant N_PF_IP_CORE_OUT_CHANS : natural := 42;
  --constant N_CHANS_PER_CORE : natural := 12;
  --constant PF_RESHAPE_FACTOR : natural := 6;
  
  constant N_IN_CHANS  : natural := 42;
  constant N_OUT_CHANS : natural := 42;
  
end;
    
