library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library IO;
use IO.DataType.all;
use IO.ArrayTypes.all;

library JetCompute;

use work.PkgConstants.all;

entity JetComputeWrapped is
port(
    clk : in std_logic;
    sum_pts : in Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    sum_pt_etas : in Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    sum_pt_phis : in Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    seed_eta : in tData := cNull;
    seed_phi : in tData := cNull;
    jet : out tData := cNull
);
end JetComputeWrapped;

architecture rtl of JetComputeWrapped is
    signal jeti : tData := cNull;
begin

    HLSIP : entity JetCompute.jet_compute
    port map(
    ap_clk => clk,
    ap_rst => '0',
    ap_start => '1',
    sum_pts_0_V => sum_pts(0).data(15 downto 0),
    sum_pts_1_V => sum_pts(1).data(15 downto 0),
    sum_pts_2_V => sum_pts(2).data(15 downto 0),
    sum_pts_3_V => sum_pts(3).data(15 downto 0),
    sum_pts_4_V => sum_pts(4).data(15 downto 0),
    sum_pts_5_V => sum_pts(5).data(15 downto 0),
    sum_pts_6_V => sum_pts(6).data(15 downto 0),
    sum_pts_7_V => sum_pts(7).data(15 downto 0),
    sum_pts_8_V => sum_pts(8).data(15 downto 0),
    sum_pts_9_V => sum_pts(9).data(15 downto 0),
    sum_pts_10_V => sum_pts(10).data(15 downto 0),
    sum_pts_11_V => sum_pts(11).data(15 downto 0),
    sum_pts_12_V => sum_pts(12).data(15 downto 0),
    sum_pts_13_V => sum_pts(13).data(15 downto 0),
    sum_pts_14_V => sum_pts(14).data(15 downto 0),
    sum_pts_15_V => sum_pts(15).data(15 downto 0),
    sum_pts_16_V => sum_pts(16).data(15 downto 0),
    sum_pts_17_V => sum_pts(17).data(15 downto 0),
    sum_pts_18_V => sum_pts(18).data(15 downto 0),
    sum_pts_19_V => sum_pts(19).data(15 downto 0),
    sum_pts_20_V => sum_pts(20).data(15 downto 0),
    sum_pts_21_V => sum_pts(21).data(15 downto 0),
    sum_pts_22_V => sum_pts(22).data(15 downto 0),
    sum_pts_23_V => sum_pts(23).data(15 downto 0),
    sum_pts_24_V => sum_pts(24).data(15 downto 0),
    sum_pts_25_V => sum_pts(25).data(15 downto 0),
    sum_pts_26_V => sum_pts(26).data(15 downto 0),
    sum_pts_27_V => sum_pts(27).data(15 downto 0),
    sum_pts_28_V => sum_pts(28).data(15 downto 0),
    sum_pts_29_V => sum_pts(29).data(15 downto 0),
    sum_pts_30_V => sum_pts(30).data(15 downto 0),
    sum_pts_31_V => sum_pts(31).data(15 downto 0),
    sum_pts_32_V => sum_pts(32).data(15 downto 0),
    sum_pts_33_V => sum_pts(33).data(15 downto 0),
    sum_pts_34_V => sum_pts(34).data(15 downto 0),
    sum_pts_35_V => sum_pts(35).data(15 downto 0),
    sum_pts_36_V => sum_pts(36).data(15 downto 0),
    sum_pts_37_V => sum_pts(37).data(15 downto 0),
    sum_pts_38_V => sum_pts(38).data(15 downto 0),
    sum_pts_39_V => sum_pts(39).data(15 downto 0),
    sum_pts_40_V => sum_pts(40).data(15 downto 0),
    sum_pts_41_V => sum_pts(41).data(15 downto 0),
    sum_pts_42_V => sum_pts(42).data(15 downto 0),
    sum_pts_43_V => sum_pts(43).data(15 downto 0),
    sum_pts_44_V => sum_pts(44).data(15 downto 0),
    sum_pts_45_V => sum_pts(45).data(15 downto 0),
    sum_pts_46_V => sum_pts(46).data(15 downto 0),
    sum_pts_47_V => sum_pts(47).data(15 downto 0),
    sum_pts_48_V => sum_pts(48).data(15 downto 0),
    sum_pts_49_V => sum_pts(49).data(15 downto 0),
    sum_pts_50_V => sum_pts(50).data(15 downto 0),
    sum_pts_51_V => sum_pts(51).data(15 downto 0),
    sum_pts_52_V => sum_pts(52).data(15 downto 0),
    sum_pts_53_V => sum_pts(53).data(15 downto 0),
    sum_pts_54_V => sum_pts(54).data(15 downto 0),
    sum_pts_55_V => sum_pts(55).data(15 downto 0),
    sum_pts_56_V => sum_pts(56).data(15 downto 0),
    sum_pts_57_V => sum_pts(57).data(15 downto 0),
    sum_pts_58_V => sum_pts(58).data(15 downto 0),
    sum_pts_59_V => sum_pts(59).data(15 downto 0),
    sum_pts_60_V => sum_pts(60).data(15 downto 0),
    sum_pts_61_V => sum_pts(61).data(15 downto 0),
    sum_pts_62_V => sum_pts(62).data(15 downto 0),
    sum_pts_63_V => sum_pts(63).data(15 downto 0),
    sum_pts_64_V => sum_pts(64).data(15 downto 0),
    sum_pts_65_V => sum_pts(65).data(15 downto 0),
    sum_pts_66_V => sum_pts(66).data(15 downto 0),
    sum_pts_67_V => sum_pts(67).data(15 downto 0),
    sum_pts_68_V => sum_pts(68).data(15 downto 0),
    sum_pts_69_V => sum_pts(69).data(15 downto 0),
    sum_pts_70_V => sum_pts(70).data(15 downto 0),
    sum_pts_71_V => sum_pts(71).data(15 downto 0),
    sum_pts_72_V => sum_pts(72).data(15 downto 0),
    sum_pts_73_V => sum_pts(73).data(15 downto 0),
    sum_pts_74_V => sum_pts(74).data(15 downto 0),
    sum_pts_75_V => sum_pts(75).data(15 downto 0),
    sum_pts_76_V => sum_pts(76).data(15 downto 0),
    sum_pts_77_V => sum_pts(77).data(15 downto 0),
    sum_pts_78_V => sum_pts(78).data(15 downto 0),
    sum_pts_79_V => sum_pts(79).data(15 downto 0),
    sum_pts_80_V => sum_pts(80).data(15 downto 0),
    sum_pts_81_V => sum_pts(81).data(15 downto 0),
    sum_pts_82_V => sum_pts(82).data(15 downto 0),
    sum_pts_83_V => sum_pts(83).data(15 downto 0),
    sum_pts_84_V => sum_pts(84).data(15 downto 0),
    sum_pts_85_V => sum_pts(85).data(15 downto 0),
    sum_pts_86_V => sum_pts(86).data(15 downto 0),
    sum_pts_87_V => sum_pts(87).data(15 downto 0),
    sum_pts_88_V => sum_pts(88).data(15 downto 0),
    sum_pts_89_V => sum_pts(89).data(15 downto 0),
    sum_pts_90_V => sum_pts(90).data(15 downto 0),
    sum_pts_91_V => sum_pts(91).data(15 downto 0),
    sum_pts_92_V => sum_pts(92).data(15 downto 0),
    sum_pts_93_V => sum_pts(93).data(15 downto 0),
    sum_pts_94_V => sum_pts(94).data(15 downto 0),
    sum_pts_95_V => sum_pts(95).data(15 downto 0),
    sum_pts_96_V => sum_pts(96).data(15 downto 0),
    sum_pts_97_V => sum_pts(97).data(15 downto 0),
    sum_pts_98_V => sum_pts(98).data(15 downto 0),
    sum_pts_99_V => sum_pts(99).data(15 downto 0),
    sum_pts_100_V => sum_pts(100).data(15 downto 0),
    sum_pts_101_V => sum_pts(101).data(15 downto 0),
    sum_pts_102_V => sum_pts(102).data(15 downto 0),
    sum_pts_103_V => sum_pts(103).data(15 downto 0),
    sum_pts_104_V => sum_pts(104).data(15 downto 0),
    sum_pts_105_V => sum_pts(105).data(15 downto 0),
    sum_pts_106_V => sum_pts(106).data(15 downto 0),
    sum_pts_107_V => sum_pts(107).data(15 downto 0),
    sum_pts_108_V => sum_pts(108).data(15 downto 0),
    sum_pts_109_V => sum_pts(109).data(15 downto 0),
    sum_pts_110_V => sum_pts(110).data(15 downto 0),
    sum_pts_111_V => sum_pts(111).data(15 downto 0),
    sum_pts_112_V => sum_pts(112).data(15 downto 0),
    sum_pts_113_V => sum_pts(113).data(15 downto 0),
    sum_pts_114_V => sum_pts(114).data(15 downto 0),
    sum_pts_115_V => sum_pts(115).data(15 downto 0),
    sum_pts_116_V => sum_pts(116).data(15 downto 0),
    sum_pts_117_V => sum_pts(117).data(15 downto 0),
    sum_pts_118_V => sum_pts(118).data(15 downto 0),
    sum_pts_119_V => sum_pts(119).data(15 downto 0),
    sum_pts_120_V => sum_pts(120).data(15 downto 0),
    sum_pts_121_V => sum_pts(121).data(15 downto 0),
    sum_pts_122_V => sum_pts(122).data(15 downto 0),
    sum_pts_123_V => sum_pts(123).data(15 downto 0),
    sum_pts_124_V => sum_pts(124).data(15 downto 0),
    sum_pts_125_V => sum_pts(125).data(15 downto 0),
    sum_pts_126_V => sum_pts(126).data(15 downto 0),
    sum_pts_127_V => sum_pts(127).data(15 downto 0),
    sum_pt_etas_0_V => sum_pt_etas(0).data(21 downto 0),
    sum_pt_etas_1_V => sum_pt_etas(1).data(21 downto 0),
    sum_pt_etas_2_V => sum_pt_etas(2).data(21 downto 0),
    sum_pt_etas_3_V => sum_pt_etas(3).data(21 downto 0),
    sum_pt_etas_4_V => sum_pt_etas(4).data(21 downto 0),
    sum_pt_etas_5_V => sum_pt_etas(5).data(21 downto 0),
    sum_pt_etas_6_V => sum_pt_etas(6).data(21 downto 0),
    sum_pt_etas_7_V => sum_pt_etas(7).data(21 downto 0),
    sum_pt_etas_8_V => sum_pt_etas(8).data(21 downto 0),
    sum_pt_etas_9_V => sum_pt_etas(9).data(21 downto 0),
    sum_pt_etas_10_V => sum_pt_etas(10).data(21 downto 0),
    sum_pt_etas_11_V => sum_pt_etas(11).data(21 downto 0),
    sum_pt_etas_12_V => sum_pt_etas(12).data(21 downto 0),
    sum_pt_etas_13_V => sum_pt_etas(13).data(21 downto 0),
    sum_pt_etas_14_V => sum_pt_etas(14).data(21 downto 0),
    sum_pt_etas_15_V => sum_pt_etas(15).data(21 downto 0),
    sum_pt_etas_16_V => sum_pt_etas(16).data(21 downto 0),
    sum_pt_etas_17_V => sum_pt_etas(17).data(21 downto 0),
    sum_pt_etas_18_V => sum_pt_etas(18).data(21 downto 0),
    sum_pt_etas_19_V => sum_pt_etas(19).data(21 downto 0),
    sum_pt_etas_20_V => sum_pt_etas(20).data(21 downto 0),
    sum_pt_etas_21_V => sum_pt_etas(21).data(21 downto 0),
    sum_pt_etas_22_V => sum_pt_etas(22).data(21 downto 0),
    sum_pt_etas_23_V => sum_pt_etas(23).data(21 downto 0),
    sum_pt_etas_24_V => sum_pt_etas(24).data(21 downto 0),
    sum_pt_etas_25_V => sum_pt_etas(25).data(21 downto 0),
    sum_pt_etas_26_V => sum_pt_etas(26).data(21 downto 0),
    sum_pt_etas_27_V => sum_pt_etas(27).data(21 downto 0),
    sum_pt_etas_28_V => sum_pt_etas(28).data(21 downto 0),
    sum_pt_etas_29_V => sum_pt_etas(29).data(21 downto 0),
    sum_pt_etas_30_V => sum_pt_etas(30).data(21 downto 0),
    sum_pt_etas_31_V => sum_pt_etas(31).data(21 downto 0),
    sum_pt_etas_32_V => sum_pt_etas(32).data(21 downto 0),
    sum_pt_etas_33_V => sum_pt_etas(33).data(21 downto 0),
    sum_pt_etas_34_V => sum_pt_etas(34).data(21 downto 0),
    sum_pt_etas_35_V => sum_pt_etas(35).data(21 downto 0),
    sum_pt_etas_36_V => sum_pt_etas(36).data(21 downto 0),
    sum_pt_etas_37_V => sum_pt_etas(37).data(21 downto 0),
    sum_pt_etas_38_V => sum_pt_etas(38).data(21 downto 0),
    sum_pt_etas_39_V => sum_pt_etas(39).data(21 downto 0),
    sum_pt_etas_40_V => sum_pt_etas(40).data(21 downto 0),
    sum_pt_etas_41_V => sum_pt_etas(41).data(21 downto 0),
    sum_pt_etas_42_V => sum_pt_etas(42).data(21 downto 0),
    sum_pt_etas_43_V => sum_pt_etas(43).data(21 downto 0),
    sum_pt_etas_44_V => sum_pt_etas(44).data(21 downto 0),
    sum_pt_etas_45_V => sum_pt_etas(45).data(21 downto 0),
    sum_pt_etas_46_V => sum_pt_etas(46).data(21 downto 0),
    sum_pt_etas_47_V => sum_pt_etas(47).data(21 downto 0),
    sum_pt_etas_48_V => sum_pt_etas(48).data(21 downto 0),
    sum_pt_etas_49_V => sum_pt_etas(49).data(21 downto 0),
    sum_pt_etas_50_V => sum_pt_etas(50).data(21 downto 0),
    sum_pt_etas_51_V => sum_pt_etas(51).data(21 downto 0),
    sum_pt_etas_52_V => sum_pt_etas(52).data(21 downto 0),
    sum_pt_etas_53_V => sum_pt_etas(53).data(21 downto 0),
    sum_pt_etas_54_V => sum_pt_etas(54).data(21 downto 0),
    sum_pt_etas_55_V => sum_pt_etas(55).data(21 downto 0),
    sum_pt_etas_56_V => sum_pt_etas(56).data(21 downto 0),
    sum_pt_etas_57_V => sum_pt_etas(57).data(21 downto 0),
    sum_pt_etas_58_V => sum_pt_etas(58).data(21 downto 0),
    sum_pt_etas_59_V => sum_pt_etas(59).data(21 downto 0),
    sum_pt_etas_60_V => sum_pt_etas(60).data(21 downto 0),
    sum_pt_etas_61_V => sum_pt_etas(61).data(21 downto 0),
    sum_pt_etas_62_V => sum_pt_etas(62).data(21 downto 0),
    sum_pt_etas_63_V => sum_pt_etas(63).data(21 downto 0),
    sum_pt_etas_64_V => sum_pt_etas(64).data(21 downto 0),
    sum_pt_etas_65_V => sum_pt_etas(65).data(21 downto 0),
    sum_pt_etas_66_V => sum_pt_etas(66).data(21 downto 0),
    sum_pt_etas_67_V => sum_pt_etas(67).data(21 downto 0),
    sum_pt_etas_68_V => sum_pt_etas(68).data(21 downto 0),
    sum_pt_etas_69_V => sum_pt_etas(69).data(21 downto 0),
    sum_pt_etas_70_V => sum_pt_etas(70).data(21 downto 0),
    sum_pt_etas_71_V => sum_pt_etas(71).data(21 downto 0),
    sum_pt_etas_72_V => sum_pt_etas(72).data(21 downto 0),
    sum_pt_etas_73_V => sum_pt_etas(73).data(21 downto 0),
    sum_pt_etas_74_V => sum_pt_etas(74).data(21 downto 0),
    sum_pt_etas_75_V => sum_pt_etas(75).data(21 downto 0),
    sum_pt_etas_76_V => sum_pt_etas(76).data(21 downto 0),
    sum_pt_etas_77_V => sum_pt_etas(77).data(21 downto 0),
    sum_pt_etas_78_V => sum_pt_etas(78).data(21 downto 0),
    sum_pt_etas_79_V => sum_pt_etas(79).data(21 downto 0),
    sum_pt_etas_80_V => sum_pt_etas(80).data(21 downto 0),
    sum_pt_etas_81_V => sum_pt_etas(81).data(21 downto 0),
    sum_pt_etas_82_V => sum_pt_etas(82).data(21 downto 0),
    sum_pt_etas_83_V => sum_pt_etas(83).data(21 downto 0),
    sum_pt_etas_84_V => sum_pt_etas(84).data(21 downto 0),
    sum_pt_etas_85_V => sum_pt_etas(85).data(21 downto 0),
    sum_pt_etas_86_V => sum_pt_etas(86).data(21 downto 0),
    sum_pt_etas_87_V => sum_pt_etas(87).data(21 downto 0),
    sum_pt_etas_88_V => sum_pt_etas(88).data(21 downto 0),
    sum_pt_etas_89_V => sum_pt_etas(89).data(21 downto 0),
    sum_pt_etas_90_V => sum_pt_etas(90).data(21 downto 0),
    sum_pt_etas_91_V => sum_pt_etas(91).data(21 downto 0),
    sum_pt_etas_92_V => sum_pt_etas(92).data(21 downto 0),
    sum_pt_etas_93_V => sum_pt_etas(93).data(21 downto 0),
    sum_pt_etas_94_V => sum_pt_etas(94).data(21 downto 0),
    sum_pt_etas_95_V => sum_pt_etas(95).data(21 downto 0),
    sum_pt_etas_96_V => sum_pt_etas(96).data(21 downto 0),
    sum_pt_etas_97_V => sum_pt_etas(97).data(21 downto 0),
    sum_pt_etas_98_V => sum_pt_etas(98).data(21 downto 0),
    sum_pt_etas_99_V => sum_pt_etas(99).data(21 downto 0),
    sum_pt_etas_100_V => sum_pt_etas(100).data(21 downto 0),
    sum_pt_etas_101_V => sum_pt_etas(101).data(21 downto 0),
    sum_pt_etas_102_V => sum_pt_etas(102).data(21 downto 0),
    sum_pt_etas_103_V => sum_pt_etas(103).data(21 downto 0),
    sum_pt_etas_104_V => sum_pt_etas(104).data(21 downto 0),
    sum_pt_etas_105_V => sum_pt_etas(105).data(21 downto 0),
    sum_pt_etas_106_V => sum_pt_etas(106).data(21 downto 0),
    sum_pt_etas_107_V => sum_pt_etas(107).data(21 downto 0),
    sum_pt_etas_108_V => sum_pt_etas(108).data(21 downto 0),
    sum_pt_etas_109_V => sum_pt_etas(109).data(21 downto 0),
    sum_pt_etas_110_V => sum_pt_etas(110).data(21 downto 0),
    sum_pt_etas_111_V => sum_pt_etas(111).data(21 downto 0),
    sum_pt_etas_112_V => sum_pt_etas(112).data(21 downto 0),
    sum_pt_etas_113_V => sum_pt_etas(113).data(21 downto 0),
    sum_pt_etas_114_V => sum_pt_etas(114).data(21 downto 0),
    sum_pt_etas_115_V => sum_pt_etas(115).data(21 downto 0),
    sum_pt_etas_116_V => sum_pt_etas(116).data(21 downto 0),
    sum_pt_etas_117_V => sum_pt_etas(117).data(21 downto 0),
    sum_pt_etas_118_V => sum_pt_etas(118).data(21 downto 0),
    sum_pt_etas_119_V => sum_pt_etas(119).data(21 downto 0),
    sum_pt_etas_120_V => sum_pt_etas(120).data(21 downto 0),
    sum_pt_etas_121_V => sum_pt_etas(121).data(21 downto 0),
    sum_pt_etas_122_V => sum_pt_etas(122).data(21 downto 0),
    sum_pt_etas_123_V => sum_pt_etas(123).data(21 downto 0),
    sum_pt_etas_124_V => sum_pt_etas(124).data(21 downto 0),
    sum_pt_etas_125_V => sum_pt_etas(125).data(21 downto 0),
    sum_pt_etas_126_V => sum_pt_etas(126).data(21 downto 0),
    sum_pt_etas_127_V => sum_pt_etas(127).data(21 downto 0),
    sum_pt_phis_0_V => sum_pt_phis(0).data(21 downto 0),
    sum_pt_phis_1_V => sum_pt_phis(1).data(21 downto 0),
    sum_pt_phis_2_V => sum_pt_phis(2).data(21 downto 0),
    sum_pt_phis_3_V => sum_pt_phis(3).data(21 downto 0),
    sum_pt_phis_4_V => sum_pt_phis(4).data(21 downto 0),
    sum_pt_phis_5_V => sum_pt_phis(5).data(21 downto 0),
    sum_pt_phis_6_V => sum_pt_phis(6).data(21 downto 0),
    sum_pt_phis_7_V => sum_pt_phis(7).data(21 downto 0),
    sum_pt_phis_8_V => sum_pt_phis(8).data(21 downto 0),
    sum_pt_phis_9_V => sum_pt_phis(9).data(21 downto 0),
    sum_pt_phis_10_V => sum_pt_phis(10).data(21 downto 0),
    sum_pt_phis_11_V => sum_pt_phis(11).data(21 downto 0),
    sum_pt_phis_12_V => sum_pt_phis(12).data(21 downto 0),
    sum_pt_phis_13_V => sum_pt_phis(13).data(21 downto 0),
    sum_pt_phis_14_V => sum_pt_phis(14).data(21 downto 0),
    sum_pt_phis_15_V => sum_pt_phis(15).data(21 downto 0),
    sum_pt_phis_16_V => sum_pt_phis(16).data(21 downto 0),
    sum_pt_phis_17_V => sum_pt_phis(17).data(21 downto 0),
    sum_pt_phis_18_V => sum_pt_phis(18).data(21 downto 0),
    sum_pt_phis_19_V => sum_pt_phis(19).data(21 downto 0),
    sum_pt_phis_20_V => sum_pt_phis(20).data(21 downto 0),
    sum_pt_phis_21_V => sum_pt_phis(21).data(21 downto 0),
    sum_pt_phis_22_V => sum_pt_phis(22).data(21 downto 0),
    sum_pt_phis_23_V => sum_pt_phis(23).data(21 downto 0),
    sum_pt_phis_24_V => sum_pt_phis(24).data(21 downto 0),
    sum_pt_phis_25_V => sum_pt_phis(25).data(21 downto 0),
    sum_pt_phis_26_V => sum_pt_phis(26).data(21 downto 0),
    sum_pt_phis_27_V => sum_pt_phis(27).data(21 downto 0),
    sum_pt_phis_28_V => sum_pt_phis(28).data(21 downto 0),
    sum_pt_phis_29_V => sum_pt_phis(29).data(21 downto 0),
    sum_pt_phis_30_V => sum_pt_phis(30).data(21 downto 0),
    sum_pt_phis_31_V => sum_pt_phis(31).data(21 downto 0),
    sum_pt_phis_32_V => sum_pt_phis(32).data(21 downto 0),
    sum_pt_phis_33_V => sum_pt_phis(33).data(21 downto 0),
    sum_pt_phis_34_V => sum_pt_phis(34).data(21 downto 0),
    sum_pt_phis_35_V => sum_pt_phis(35).data(21 downto 0),
    sum_pt_phis_36_V => sum_pt_phis(36).data(21 downto 0),
    sum_pt_phis_37_V => sum_pt_phis(37).data(21 downto 0),
    sum_pt_phis_38_V => sum_pt_phis(38).data(21 downto 0),
    sum_pt_phis_39_V => sum_pt_phis(39).data(21 downto 0),
    sum_pt_phis_40_V => sum_pt_phis(40).data(21 downto 0),
    sum_pt_phis_41_V => sum_pt_phis(41).data(21 downto 0),
    sum_pt_phis_42_V => sum_pt_phis(42).data(21 downto 0),
    sum_pt_phis_43_V => sum_pt_phis(43).data(21 downto 0),
    sum_pt_phis_44_V => sum_pt_phis(44).data(21 downto 0),
    sum_pt_phis_45_V => sum_pt_phis(45).data(21 downto 0),
    sum_pt_phis_46_V => sum_pt_phis(46).data(21 downto 0),
    sum_pt_phis_47_V => sum_pt_phis(47).data(21 downto 0),
    sum_pt_phis_48_V => sum_pt_phis(48).data(21 downto 0),
    sum_pt_phis_49_V => sum_pt_phis(49).data(21 downto 0),
    sum_pt_phis_50_V => sum_pt_phis(50).data(21 downto 0),
    sum_pt_phis_51_V => sum_pt_phis(51).data(21 downto 0),
    sum_pt_phis_52_V => sum_pt_phis(52).data(21 downto 0),
    sum_pt_phis_53_V => sum_pt_phis(53).data(21 downto 0),
    sum_pt_phis_54_V => sum_pt_phis(54).data(21 downto 0),
    sum_pt_phis_55_V => sum_pt_phis(55).data(21 downto 0),
    sum_pt_phis_56_V => sum_pt_phis(56).data(21 downto 0),
    sum_pt_phis_57_V => sum_pt_phis(57).data(21 downto 0),
    sum_pt_phis_58_V => sum_pt_phis(58).data(21 downto 0),
    sum_pt_phis_59_V => sum_pt_phis(59).data(21 downto 0),
    sum_pt_phis_60_V => sum_pt_phis(60).data(21 downto 0),
    sum_pt_phis_61_V => sum_pt_phis(61).data(21 downto 0),
    sum_pt_phis_62_V => sum_pt_phis(62).data(21 downto 0),
    sum_pt_phis_63_V => sum_pt_phis(63).data(21 downto 0),
    sum_pt_phis_64_V => sum_pt_phis(64).data(21 downto 0),
    sum_pt_phis_65_V => sum_pt_phis(65).data(21 downto 0),
    sum_pt_phis_66_V => sum_pt_phis(66).data(21 downto 0),
    sum_pt_phis_67_V => sum_pt_phis(67).data(21 downto 0),
    sum_pt_phis_68_V => sum_pt_phis(68).data(21 downto 0),
    sum_pt_phis_69_V => sum_pt_phis(69).data(21 downto 0),
    sum_pt_phis_70_V => sum_pt_phis(70).data(21 downto 0),
    sum_pt_phis_71_V => sum_pt_phis(71).data(21 downto 0),
    sum_pt_phis_72_V => sum_pt_phis(72).data(21 downto 0),
    sum_pt_phis_73_V => sum_pt_phis(73).data(21 downto 0),
    sum_pt_phis_74_V => sum_pt_phis(74).data(21 downto 0),
    sum_pt_phis_75_V => sum_pt_phis(75).data(21 downto 0),
    sum_pt_phis_76_V => sum_pt_phis(76).data(21 downto 0),
    sum_pt_phis_77_V => sum_pt_phis(77).data(21 downto 0),
    sum_pt_phis_78_V => sum_pt_phis(78).data(21 downto 0),
    sum_pt_phis_79_V => sum_pt_phis(79).data(21 downto 0),
    sum_pt_phis_80_V => sum_pt_phis(80).data(21 downto 0),
    sum_pt_phis_81_V => sum_pt_phis(81).data(21 downto 0),
    sum_pt_phis_82_V => sum_pt_phis(82).data(21 downto 0),
    sum_pt_phis_83_V => sum_pt_phis(83).data(21 downto 0),
    sum_pt_phis_84_V => sum_pt_phis(84).data(21 downto 0),
    sum_pt_phis_85_V => sum_pt_phis(85).data(21 downto 0),
    sum_pt_phis_86_V => sum_pt_phis(86).data(21 downto 0),
    sum_pt_phis_87_V => sum_pt_phis(87).data(21 downto 0),
    sum_pt_phis_88_V => sum_pt_phis(88).data(21 downto 0),
    sum_pt_phis_89_V => sum_pt_phis(89).data(21 downto 0),
    sum_pt_phis_90_V => sum_pt_phis(90).data(21 downto 0),
    sum_pt_phis_91_V => sum_pt_phis(91).data(21 downto 0),
    sum_pt_phis_92_V => sum_pt_phis(92).data(21 downto 0),
    sum_pt_phis_93_V => sum_pt_phis(93).data(21 downto 0),
    sum_pt_phis_94_V => sum_pt_phis(94).data(21 downto 0),
    sum_pt_phis_95_V => sum_pt_phis(95).data(21 downto 0),
    sum_pt_phis_96_V => sum_pt_phis(96).data(21 downto 0),
    sum_pt_phis_97_V => sum_pt_phis(97).data(21 downto 0),
    sum_pt_phis_98_V => sum_pt_phis(98).data(21 downto 0),
    sum_pt_phis_99_V => sum_pt_phis(99).data(21 downto 0),
    sum_pt_phis_100_V => sum_pt_phis(100).data(21 downto 0),
    sum_pt_phis_101_V => sum_pt_phis(101).data(21 downto 0),
    sum_pt_phis_102_V => sum_pt_phis(102).data(21 downto 0),
    sum_pt_phis_103_V => sum_pt_phis(103).data(21 downto 0),
    sum_pt_phis_104_V => sum_pt_phis(104).data(21 downto 0),
    sum_pt_phis_105_V => sum_pt_phis(105).data(21 downto 0),
    sum_pt_phis_106_V => sum_pt_phis(106).data(21 downto 0),
    sum_pt_phis_107_V => sum_pt_phis(107).data(21 downto 0),
    sum_pt_phis_108_V => sum_pt_phis(108).data(21 downto 0),
    sum_pt_phis_109_V => sum_pt_phis(109).data(21 downto 0),
    sum_pt_phis_110_V => sum_pt_phis(110).data(21 downto 0),
    sum_pt_phis_111_V => sum_pt_phis(111).data(21 downto 0),
    sum_pt_phis_112_V => sum_pt_phis(112).data(21 downto 0),
    sum_pt_phis_113_V => sum_pt_phis(113).data(21 downto 0),
    sum_pt_phis_114_V => sum_pt_phis(114).data(21 downto 0),
    sum_pt_phis_115_V => sum_pt_phis(115).data(21 downto 0),
    sum_pt_phis_116_V => sum_pt_phis(116).data(21 downto 0),
    sum_pt_phis_117_V => sum_pt_phis(117).data(21 downto 0),
    sum_pt_phis_118_V => sum_pt_phis(118).data(21 downto 0),
    sum_pt_phis_119_V => sum_pt_phis(119).data(21 downto 0),
    sum_pt_phis_120_V => sum_pt_phis(120).data(21 downto 0),
    sum_pt_phis_121_V => sum_pt_phis(121).data(21 downto 0),
    sum_pt_phis_122_V => sum_pt_phis(122).data(21 downto 0),
    sum_pt_phis_123_V => sum_pt_phis(123).data(21 downto 0),
    sum_pt_phis_124_V => sum_pt_phis(124).data(21 downto 0),
    sum_pt_phis_125_V => sum_pt_phis(125).data(21 downto 0),
    sum_pt_phis_126_V => sum_pt_phis(126).data(21 downto 0),
    sum_pt_phis_127_V => sum_pt_phis(127).data(21 downto 0),
    seed_eta_V => seed_eta.data(9 downto 0),
    seed_phi_V => seed_phi.data(9 downto 0),
    jet => jet.data(45 downto 0)
    );

end rtl;
