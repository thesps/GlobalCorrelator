../../../../../../RuflCore/firmware/hdl/ReuseableElements/PairReduceMax.vhd