../../../../../../../GlobalCorrelator_HLS/JetLoop/solution1/syn/vhdl/jet_loop_mul_mul_dEe.vhd