../../../../../../../GlobalCorrelator_HLS/JetLoop/solution1/syn/vhdl/dreg_ap_fixed_s.vhd