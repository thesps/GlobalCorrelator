library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library IO;
use IO.DataType.all;
use IO.ArrayTypes.all;

library JetLoop;

use work.PkgConstants.all;

entity JetLoopWrapped is
port(
    clk : in std_logic;
    particles_in : in Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    particles_out : out Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    partialParts : out Vector(0 to NPARTICLES-1) := NullVector(NPARTICLES);
    seed_eta : out tData := cNull;
    seed_phi : out tData := cNull
);
end JetLoopWrapped;

architecture rtl of JetLoopWrapped is

begin

    HLSIP : entity JetLoop.jet_loop
    port map(
    ap_clk => clk,
    ap_rst => '0',
    ap_start => '1',
    particles_in_0 => particles_in(0).data(35 downto 0),
    particles_in_1 => particles_in(1).data(35 downto 0),
    particles_in_2 => particles_in(2).data(35 downto 0),
    particles_in_3 => particles_in(3).data(35 downto 0),
    particles_in_4 => particles_in(4).data(35 downto 0),
    particles_in_5 => particles_in(5).data(35 downto 0),
    particles_in_6 => particles_in(6).data(35 downto 0),
    particles_in_7 => particles_in(7).data(35 downto 0),
    particles_in_8 => particles_in(8).data(35 downto 0),
    particles_in_9 => particles_in(9).data(35 downto 0),
    particles_in_10 => particles_in(10).data(35 downto 0),
    particles_in_11 => particles_in(11).data(35 downto 0),
    particles_in_12 => particles_in(12).data(35 downto 0),
    particles_in_13 => particles_in(13).data(35 downto 0),
    particles_in_14 => particles_in(14).data(35 downto 0),
    particles_in_15 => particles_in(15).data(35 downto 0),
    particles_in_16 => particles_in(16).data(35 downto 0),
    particles_in_17 => particles_in(17).data(35 downto 0),
    particles_in_18 => particles_in(18).data(35 downto 0),
    particles_in_19 => particles_in(19).data(35 downto 0),
    particles_in_20 => particles_in(20).data(35 downto 0),
    particles_in_21 => particles_in(21).data(35 downto 0),
    particles_in_22 => particles_in(22).data(35 downto 0),
    particles_in_23 => particles_in(23).data(35 downto 0),
    particles_in_24 => particles_in(24).data(35 downto 0),
    particles_in_25 => particles_in(25).data(35 downto 0),
    particles_in_26 => particles_in(26).data(35 downto 0),
    particles_in_27 => particles_in(27).data(35 downto 0),
    particles_in_28 => particles_in(28).data(35 downto 0),
    particles_in_29 => particles_in(29).data(35 downto 0),
    particles_in_30 => particles_in(30).data(35 downto 0),
    particles_in_31 => particles_in(31).data(35 downto 0),
    particles_in_32 => particles_in(32).data(35 downto 0),
    particles_in_33 => particles_in(33).data(35 downto 0),
    particles_in_34 => particles_in(34).data(35 downto 0),
    particles_in_35 => particles_in(35).data(35 downto 0),
    particles_in_36 => particles_in(36).data(35 downto 0),
    particles_in_37 => particles_in(37).data(35 downto 0),
    particles_in_38 => particles_in(38).data(35 downto 0),
    particles_in_39 => particles_in(39).data(35 downto 0),
    particles_in_40 => particles_in(40).data(35 downto 0),
    particles_in_41 => particles_in(41).data(35 downto 0),
    particles_in_42 => particles_in(42).data(35 downto 0),
    particles_in_43 => particles_in(43).data(35 downto 0),
    particles_in_44 => particles_in(44).data(35 downto 0),
    particles_in_45 => particles_in(45).data(35 downto 0),
    particles_in_46 => particles_in(46).data(35 downto 0),
    particles_in_47 => particles_in(47).data(35 downto 0),
    particles_in_48 => particles_in(48).data(35 downto 0),
    particles_in_49 => particles_in(49).data(35 downto 0),
    particles_in_50 => particles_in(50).data(35 downto 0),
    particles_in_51 => particles_in(51).data(35 downto 0),
    particles_in_52 => particles_in(52).data(35 downto 0),
    particles_in_53 => particles_in(53).data(35 downto 0),
    particles_in_54 => particles_in(54).data(35 downto 0),
    particles_in_55 => particles_in(55).data(35 downto 0),
    particles_in_56 => particles_in(56).data(35 downto 0),
    particles_in_57 => particles_in(57).data(35 downto 0),
    particles_in_58 => particles_in(58).data(35 downto 0),
    particles_in_59 => particles_in(59).data(35 downto 0),
    particles_in_60 => particles_in(60).data(35 downto 0),
    particles_in_61 => particles_in(61).data(35 downto 0),
    particles_in_62 => particles_in(62).data(35 downto 0),
    particles_in_63 => particles_in(63).data(35 downto 0),
    particles_in_64 => particles_in(64).data(35 downto 0),
    particles_in_65 => particles_in(65).data(35 downto 0),
    particles_in_66 => particles_in(66).data(35 downto 0),
    particles_in_67 => particles_in(67).data(35 downto 0),
    particles_in_68 => particles_in(68).data(35 downto 0),
    particles_in_69 => particles_in(69).data(35 downto 0),
    particles_in_70 => particles_in(70).data(35 downto 0),
    particles_in_71 => particles_in(71).data(35 downto 0),
    particles_in_72 => particles_in(72).data(35 downto 0),
    particles_in_73 => particles_in(73).data(35 downto 0),
    particles_in_74 => particles_in(74).data(35 downto 0),
    particles_in_75 => particles_in(75).data(35 downto 0),
    particles_in_76 => particles_in(76).data(35 downto 0),
    particles_in_77 => particles_in(77).data(35 downto 0),
    particles_in_78 => particles_in(78).data(35 downto 0),
    particles_in_79 => particles_in(79).data(35 downto 0),
    particles_in_80 => particles_in(80).data(35 downto 0),
    particles_in_81 => particles_in(81).data(35 downto 0),
    particles_in_82 => particles_in(82).data(35 downto 0),
    particles_in_83 => particles_in(83).data(35 downto 0),
    particles_in_84 => particles_in(84).data(35 downto 0),
    particles_in_85 => particles_in(85).data(35 downto 0),
    particles_in_86 => particles_in(86).data(35 downto 0),
    particles_in_87 => particles_in(87).data(35 downto 0),
    particles_in_88 => particles_in(88).data(35 downto 0),
    particles_in_89 => particles_in(89).data(35 downto 0),
    particles_in_90 => particles_in(90).data(35 downto 0),
    particles_in_91 => particles_in(91).data(35 downto 0),
    particles_in_92 => particles_in(92).data(35 downto 0),
    particles_in_93 => particles_in(93).data(35 downto 0),
    particles_in_94 => particles_in(94).data(35 downto 0),
    particles_in_95 => particles_in(95).data(35 downto 0),
    particles_in_96 => particles_in(96).data(35 downto 0),
    particles_in_97 => particles_in(97).data(35 downto 0),
    particles_in_98 => particles_in(98).data(35 downto 0),
    particles_in_99 => particles_in(99).data(35 downto 0),
    particles_in_100 => particles_in(100).data(35 downto 0),
    particles_in_101 => particles_in(101).data(35 downto 0),
    particles_in_102 => particles_in(102).data(35 downto 0),
    particles_in_103 => particles_in(103).data(35 downto 0),
    particles_in_104 => particles_in(104).data(35 downto 0),
    particles_in_105 => particles_in(105).data(35 downto 0),
    particles_in_106 => particles_in(106).data(35 downto 0),
    particles_in_107 => particles_in(107).data(35 downto 0),
    particles_in_108 => particles_in(108).data(35 downto 0),
    particles_in_109 => particles_in(109).data(35 downto 0),
    particles_in_110 => particles_in(110).data(35 downto 0),
    particles_in_111 => particles_in(111).data(35 downto 0),
    particles_in_112 => particles_in(112).data(35 downto 0),
    particles_in_113 => particles_in(113).data(35 downto 0),
    particles_in_114 => particles_in(114).data(35 downto 0),
    particles_in_115 => particles_in(115).data(35 downto 0),
    particles_in_116 => particles_in(116).data(35 downto 0),
    particles_in_117 => particles_in(117).data(35 downto 0),
    particles_in_118 => particles_in(118).data(35 downto 0),
    particles_in_119 => particles_in(119).data(35 downto 0),
    particles_in_120 => particles_in(120).data(35 downto 0),
    particles_in_121 => particles_in(121).data(35 downto 0),
    particles_in_122 => particles_in(122).data(35 downto 0),
    particles_in_123 => particles_in(123).data(35 downto 0),
    particles_in_124 => particles_in(124).data(35 downto 0),
    particles_in_125 => particles_in(125).data(35 downto 0),
    particles_in_126 => particles_in(126).data(35 downto 0),
    particles_in_127 => particles_in(127).data(35 downto 0),
    particles_out_0 => particles_out(0).data(35 downto 0),
    particles_out_1 => particles_out(1).data(35 downto 0),
    particles_out_2 => particles_out(2).data(35 downto 0),
    particles_out_3 => particles_out(3).data(35 downto 0),
    particles_out_4 => particles_out(4).data(35 downto 0),
    particles_out_5 => particles_out(5).data(35 downto 0),
    particles_out_6 => particles_out(6).data(35 downto 0),
    particles_out_7 => particles_out(7).data(35 downto 0),
    particles_out_8 => particles_out(8).data(35 downto 0),
    particles_out_9 => particles_out(9).data(35 downto 0),
    particles_out_10 => particles_out(10).data(35 downto 0),
    particles_out_11 => particles_out(11).data(35 downto 0),
    particles_out_12 => particles_out(12).data(35 downto 0),
    particles_out_13 => particles_out(13).data(35 downto 0),
    particles_out_14 => particles_out(14).data(35 downto 0),
    particles_out_15 => particles_out(15).data(35 downto 0),
    particles_out_16 => particles_out(16).data(35 downto 0),
    particles_out_17 => particles_out(17).data(35 downto 0),
    particles_out_18 => particles_out(18).data(35 downto 0),
    particles_out_19 => particles_out(19).data(35 downto 0),
    particles_out_20 => particles_out(20).data(35 downto 0),
    particles_out_21 => particles_out(21).data(35 downto 0),
    particles_out_22 => particles_out(22).data(35 downto 0),
    particles_out_23 => particles_out(23).data(35 downto 0),
    particles_out_24 => particles_out(24).data(35 downto 0),
    particles_out_25 => particles_out(25).data(35 downto 0),
    particles_out_26 => particles_out(26).data(35 downto 0),
    particles_out_27 => particles_out(27).data(35 downto 0),
    particles_out_28 => particles_out(28).data(35 downto 0),
    particles_out_29 => particles_out(29).data(35 downto 0),
    particles_out_30 => particles_out(30).data(35 downto 0),
    particles_out_31 => particles_out(31).data(35 downto 0),
    particles_out_32 => particles_out(32).data(35 downto 0),
    particles_out_33 => particles_out(33).data(35 downto 0),
    particles_out_34 => particles_out(34).data(35 downto 0),
    particles_out_35 => particles_out(35).data(35 downto 0),
    particles_out_36 => particles_out(36).data(35 downto 0),
    particles_out_37 => particles_out(37).data(35 downto 0),
    particles_out_38 => particles_out(38).data(35 downto 0),
    particles_out_39 => particles_out(39).data(35 downto 0),
    particles_out_40 => particles_out(40).data(35 downto 0),
    particles_out_41 => particles_out(41).data(35 downto 0),
    particles_out_42 => particles_out(42).data(35 downto 0),
    particles_out_43 => particles_out(43).data(35 downto 0),
    particles_out_44 => particles_out(44).data(35 downto 0),
    particles_out_45 => particles_out(45).data(35 downto 0),
    particles_out_46 => particles_out(46).data(35 downto 0),
    particles_out_47 => particles_out(47).data(35 downto 0),
    particles_out_48 => particles_out(48).data(35 downto 0),
    particles_out_49 => particles_out(49).data(35 downto 0),
    particles_out_50 => particles_out(50).data(35 downto 0),
    particles_out_51 => particles_out(51).data(35 downto 0),
    particles_out_52 => particles_out(52).data(35 downto 0),
    particles_out_53 => particles_out(53).data(35 downto 0),
    particles_out_54 => particles_out(54).data(35 downto 0),
    particles_out_55 => particles_out(55).data(35 downto 0),
    particles_out_56 => particles_out(56).data(35 downto 0),
    particles_out_57 => particles_out(57).data(35 downto 0),
    particles_out_58 => particles_out(58).data(35 downto 0),
    particles_out_59 => particles_out(59).data(35 downto 0),
    particles_out_60 => particles_out(60).data(35 downto 0),
    particles_out_61 => particles_out(61).data(35 downto 0),
    particles_out_62 => particles_out(62).data(35 downto 0),
    particles_out_63 => particles_out(63).data(35 downto 0),
    particles_out_64 => particles_out(64).data(35 downto 0),
    particles_out_65 => particles_out(65).data(35 downto 0),
    particles_out_66 => particles_out(66).data(35 downto 0),
    particles_out_67 => particles_out(67).data(35 downto 0),
    particles_out_68 => particles_out(68).data(35 downto 0),
    particles_out_69 => particles_out(69).data(35 downto 0),
    particles_out_70 => particles_out(70).data(35 downto 0),
    particles_out_71 => particles_out(71).data(35 downto 0),
    particles_out_72 => particles_out(72).data(35 downto 0),
    particles_out_73 => particles_out(73).data(35 downto 0),
    particles_out_74 => particles_out(74).data(35 downto 0),
    particles_out_75 => particles_out(75).data(35 downto 0),
    particles_out_76 => particles_out(76).data(35 downto 0),
    particles_out_77 => particles_out(77).data(35 downto 0),
    particles_out_78 => particles_out(78).data(35 downto 0),
    particles_out_79 => particles_out(79).data(35 downto 0),
    particles_out_80 => particles_out(80).data(35 downto 0),
    particles_out_81 => particles_out(81).data(35 downto 0),
    particles_out_82 => particles_out(82).data(35 downto 0),
    particles_out_83 => particles_out(83).data(35 downto 0),
    particles_out_84 => particles_out(84).data(35 downto 0),
    particles_out_85 => particles_out(85).data(35 downto 0),
    particles_out_86 => particles_out(86).data(35 downto 0),
    particles_out_87 => particles_out(87).data(35 downto 0),
    particles_out_88 => particles_out(88).data(35 downto 0),
    particles_out_89 => particles_out(89).data(35 downto 0),
    particles_out_90 => particles_out(90).data(35 downto 0),
    particles_out_91 => particles_out(91).data(35 downto 0),
    particles_out_92 => particles_out(92).data(35 downto 0),
    particles_out_93 => particles_out(93).data(35 downto 0),
    particles_out_94 => particles_out(94).data(35 downto 0),
    particles_out_95 => particles_out(95).data(35 downto 0),
    particles_out_96 => particles_out(96).data(35 downto 0),
    particles_out_97 => particles_out(97).data(35 downto 0),
    particles_out_98 => particles_out(98).data(35 downto 0),
    particles_out_99 => particles_out(99).data(35 downto 0),
    particles_out_100 => particles_out(100).data(35 downto 0),
    particles_out_101 => particles_out(101).data(35 downto 0),
    particles_out_102 => particles_out(102).data(35 downto 0),
    particles_out_103 => particles_out(103).data(35 downto 0),
    particles_out_104 => particles_out(104).data(35 downto 0),
    particles_out_105 => particles_out(105).data(35 downto 0),
    particles_out_106 => particles_out(106).data(35 downto 0),
    particles_out_107 => particles_out(107).data(35 downto 0),
    particles_out_108 => particles_out(108).data(35 downto 0),
    particles_out_109 => particles_out(109).data(35 downto 0),
    particles_out_110 => particles_out(110).data(35 downto 0),
    particles_out_111 => particles_out(111).data(35 downto 0),
    particles_out_112 => particles_out(112).data(35 downto 0),
    particles_out_113 => particles_out(113).data(35 downto 0),
    particles_out_114 => particles_out(114).data(35 downto 0),
    particles_out_115 => particles_out(115).data(35 downto 0),
    particles_out_116 => particles_out(116).data(35 downto 0),
    particles_out_117 => particles_out(117).data(35 downto 0),
    particles_out_118 => particles_out(118).data(35 downto 0),
    particles_out_119 => particles_out(119).data(35 downto 0),
    particles_out_120 => particles_out(120).data(35 downto 0),
    particles_out_121 => particles_out(121).data(35 downto 0),
    particles_out_122 => particles_out(122).data(35 downto 0),
    particles_out_123 => particles_out(123).data(35 downto 0),
    particles_out_124 => particles_out(124).data(35 downto 0),
    particles_out_125 => particles_out(125).data(35 downto 0),
    particles_out_126 => particles_out(126).data(35 downto 0),
    particles_out_127 => particles_out(127).data(35 downto 0),
    partialParts_0 => partialParts(0).data(59 downto 0),
    partialParts_1 => partialParts(1).data(59 downto 0),
    partialParts_2 => partialParts(2).data(59 downto 0),
    partialParts_3 => partialParts(3).data(59 downto 0),
    partialParts_4 => partialParts(4).data(59 downto 0),
    partialParts_5 => partialParts(5).data(59 downto 0),
    partialParts_6 => partialParts(6).data(59 downto 0),
    partialParts_7 => partialParts(7).data(59 downto 0),
    partialParts_8 => partialParts(8).data(59 downto 0),
    partialParts_9 => partialParts(9).data(59 downto 0),
    partialParts_10 => partialParts(10).data(59 downto 0),
    partialParts_11 => partialParts(11).data(59 downto 0),
    partialParts_12 => partialParts(12).data(59 downto 0),
    partialParts_13 => partialParts(13).data(59 downto 0),
    partialParts_14 => partialParts(14).data(59 downto 0),
    partialParts_15 => partialParts(15).data(59 downto 0),
    partialParts_16 => partialParts(16).data(59 downto 0),
    partialParts_17 => partialParts(17).data(59 downto 0),
    partialParts_18 => partialParts(18).data(59 downto 0),
    partialParts_19 => partialParts(19).data(59 downto 0),
    partialParts_20 => partialParts(20).data(59 downto 0),
    partialParts_21 => partialParts(21).data(59 downto 0),
    partialParts_22 => partialParts(22).data(59 downto 0),
    partialParts_23 => partialParts(23).data(59 downto 0),
    partialParts_24 => partialParts(24).data(59 downto 0),
    partialParts_25 => partialParts(25).data(59 downto 0),
    partialParts_26 => partialParts(26).data(59 downto 0),
    partialParts_27 => partialParts(27).data(59 downto 0),
    partialParts_28 => partialParts(28).data(59 downto 0),
    partialParts_29 => partialParts(29).data(59 downto 0),
    partialParts_30 => partialParts(30).data(59 downto 0),
    partialParts_31 => partialParts(31).data(59 downto 0),
    partialParts_32 => partialParts(32).data(59 downto 0),
    partialParts_33 => partialParts(33).data(59 downto 0),
    partialParts_34 => partialParts(34).data(59 downto 0),
    partialParts_35 => partialParts(35).data(59 downto 0),
    partialParts_36 => partialParts(36).data(59 downto 0),
    partialParts_37 => partialParts(37).data(59 downto 0),
    partialParts_38 => partialParts(38).data(59 downto 0),
    partialParts_39 => partialParts(39).data(59 downto 0),
    partialParts_40 => partialParts(40).data(59 downto 0),
    partialParts_41 => partialParts(41).data(59 downto 0),
    partialParts_42 => partialParts(42).data(59 downto 0),
    partialParts_43 => partialParts(43).data(59 downto 0),
    partialParts_44 => partialParts(44).data(59 downto 0),
    partialParts_45 => partialParts(45).data(59 downto 0),
    partialParts_46 => partialParts(46).data(59 downto 0),
    partialParts_47 => partialParts(47).data(59 downto 0),
    partialParts_48 => partialParts(48).data(59 downto 0),
    partialParts_49 => partialParts(49).data(59 downto 0),
    partialParts_50 => partialParts(50).data(59 downto 0),
    partialParts_51 => partialParts(51).data(59 downto 0),
    partialParts_52 => partialParts(52).data(59 downto 0),
    partialParts_53 => partialParts(53).data(59 downto 0),
    partialParts_54 => partialParts(54).data(59 downto 0),
    partialParts_55 => partialParts(55).data(59 downto 0),
    partialParts_56 => partialParts(56).data(59 downto 0),
    partialParts_57 => partialParts(57).data(59 downto 0),
    partialParts_58 => partialParts(58).data(59 downto 0),
    partialParts_59 => partialParts(59).data(59 downto 0),
    partialParts_60 => partialParts(60).data(59 downto 0),
    partialParts_61 => partialParts(61).data(59 downto 0),
    partialParts_62 => partialParts(62).data(59 downto 0),
    partialParts_63 => partialParts(63).data(59 downto 0),
    partialParts_64 => partialParts(64).data(59 downto 0),
    partialParts_65 => partialParts(65).data(59 downto 0),
    partialParts_66 => partialParts(66).data(59 downto 0),
    partialParts_67 => partialParts(67).data(59 downto 0),
    partialParts_68 => partialParts(68).data(59 downto 0),
    partialParts_69 => partialParts(69).data(59 downto 0),
    partialParts_70 => partialParts(70).data(59 downto 0),
    partialParts_71 => partialParts(71).data(59 downto 0),
    partialParts_72 => partialParts(72).data(59 downto 0),
    partialParts_73 => partialParts(73).data(59 downto 0),
    partialParts_74 => partialParts(74).data(59 downto 0),
    partialParts_75 => partialParts(75).data(59 downto 0),
    partialParts_76 => partialParts(76).data(59 downto 0),
    partialParts_77 => partialParts(77).data(59 downto 0),
    partialParts_78 => partialParts(78).data(59 downto 0),
    partialParts_79 => partialParts(79).data(59 downto 0),
    partialParts_80 => partialParts(80).data(59 downto 0),
    partialParts_81 => partialParts(81).data(59 downto 0),
    partialParts_82 => partialParts(82).data(59 downto 0),
    partialParts_83 => partialParts(83).data(59 downto 0),
    partialParts_84 => partialParts(84).data(59 downto 0),
    partialParts_85 => partialParts(85).data(59 downto 0),
    partialParts_86 => partialParts(86).data(59 downto 0),
    partialParts_87 => partialParts(87).data(59 downto 0),
    partialParts_88 => partialParts(88).data(59 downto 0),
    partialParts_89 => partialParts(89).data(59 downto 0),
    partialParts_90 => partialParts(90).data(59 downto 0),
    partialParts_91 => partialParts(91).data(59 downto 0),
    partialParts_92 => partialParts(92).data(59 downto 0),
    partialParts_93 => partialParts(93).data(59 downto 0),
    partialParts_94 => partialParts(94).data(59 downto 0),
    partialParts_95 => partialParts(95).data(59 downto 0),
    partialParts_96 => partialParts(96).data(59 downto 0),
    partialParts_97 => partialParts(97).data(59 downto 0),
    partialParts_98 => partialParts(98).data(59 downto 0),
    partialParts_99 => partialParts(99).data(59 downto 0),
    partialParts_100 => partialParts(100).data(59 downto 0),
    partialParts_101 => partialParts(101).data(59 downto 0),
    partialParts_102 => partialParts(102).data(59 downto 0),
    partialParts_103 => partialParts(103).data(59 downto 0),
    partialParts_104 => partialParts(104).data(59 downto 0),
    partialParts_105 => partialParts(105).data(59 downto 0),
    partialParts_106 => partialParts(106).data(59 downto 0),
    partialParts_107 => partialParts(107).data(59 downto 0),
    partialParts_108 => partialParts(108).data(59 downto 0),
    partialParts_109 => partialParts(109).data(59 downto 0),
    partialParts_110 => partialParts(110).data(59 downto 0),
    partialParts_111 => partialParts(111).data(59 downto 0),
    partialParts_112 => partialParts(112).data(59 downto 0),
    partialParts_113 => partialParts(113).data(59 downto 0),
    partialParts_114 => partialParts(114).data(59 downto 0),
    partialParts_115 => partialParts(115).data(59 downto 0),
    partialParts_116 => partialParts(116).data(59 downto 0),
    partialParts_117 => partialParts(117).data(59 downto 0),
    partialParts_118 => partialParts(118).data(59 downto 0),
    partialParts_119 => partialParts(119).data(59 downto 0),
    partialParts_120 => partialParts(120).data(59 downto 0),
    partialParts_121 => partialParts(121).data(59 downto 0),
    partialParts_122 => partialParts(122).data(59 downto 0),
    partialParts_123 => partialParts(123).data(59 downto 0),
    partialParts_124 => partialParts(124).data(59 downto 0),
    partialParts_125 => partialParts(125).data(59 downto 0),
    partialParts_126 => partialParts(126).data(59 downto 0),
    partialParts_127 => partialParts(127).data(59 downto 0),
    seed_eta_V => seed_eta.data(9 downto 0),
    seed_phi_V => seed_phi.data(9 downto 0)
    );

end rtl;

